
#******
# Preview export LEF
#
#	 Preview sub-version 5.10.41.500.5.122
#
# REF LIBS: CarlPadsv2 
# TECH LIB NAME: cmos065
# TECH FILE NAME: techfile.cds
#******

VERSION 5.5 ;

NAMESCASESENSITIVE ON ;

DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

SITE IOSite
    SYMMETRY Y  ;
    CLASS PAD  ;
    SIZE 50.000 BY 75.500 ;
END IOSite

MACRO PADVDD_74x50uNOTRIG
    CLASS PAD ;
    FOREIGN PADVDD_74x50uNOTRIG 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 60.000 BY 75.500 ;
    SYMMETRY R90 ;
    SITE IOSite ;
    PIN vdd
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M1 ;
        RECT  59.500 1.300 60.000 26.500 ;
        RECT  0.000 1.300 0.500 26.500 ;
        END
    END vdd
    PIN gnd
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M1 ;
        RECT  59.495 29.000 60.000 75.500 ;
        RECT  0.000 29.000 0.500 75.500 ;
        END
    END gnd
    PIN VDDC
        DIRECTION INOUT ;
        USE POWER ;
        PORT
            CLASS CORE ;
        LAYER AP ;
        RECT  32.445 71.000 55.000 74.000 ;
        RECT  5.000 71.000 27.475 74.000 ;
        END
        PORT
            CLASS CORE ;
        LAYER M7 ;
        RECT  31.000 69.665 53.000 72.000 ;
        RECT  7.000 69.665 29.000 72.000 ;
        END
    END VDDC
    OBS
        LAYER M1 ;
        RECT  2.090 1.300 57.910 27.410 ;
        RECT  2.090 1.300 57.905 75.500 ;
        LAYER M2 ;
        RECT  0.000 1.300 60.000 26.500 ;
        RECT  0.000 36.500 60.000 37.500 ;
        RECT  0.000 39.500 60.000 40.500 ;
        RECT  1.500 1.300 58.500 75.500 ;
        RECT  0.000 47.500 60.000 75.500 ;
        LAYER M3 ;
        RECT  1.500 1.500 58.500 74.000 ;
        LAYER M4 ;
        RECT  1.500 1.500 58.500 74.000 ;
        LAYER M5 ;
        RECT  1.500 1.500 58.500 74.000 ;
        RECT  2.000 1.500 58.000 75.500 ;
        LAYER M6 ;
        RECT  1.500 1.500 58.500 74.000 ;
        RECT  2.000 1.500 58.000 75.500 ;
        LAYER M7 ;
        RECT  5.500 1.300 47.500 65.965 ;
        RECT  1.500 1.500 58.500 65.965 ;
        RECT  1.500 1.500 3.300 74.000 ;
        RECT  56.700 1.500 58.500 74.000 ;
        LAYER AP ;
        RECT  1.000 1.000 59.000 65.465 ;
        RECT  1.000 1.000 2.800 66.800 ;
        RECT  5.000 0.000 55.000 66.800 ;
        RECT  57.200 1.000 59.000 66.800 ;
    END
END PADVDD_74x50uNOTRIG

MACRO PADSPACE_C_74x74u_CH
    CLASS PAD ;
    FOREIGN PADSPACE_C_74x74u_CH 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 76.000 BY 76.000 ;
    SYMMETRY R90 ;
    SITE IOSite ;
    PIN vdd
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M1 ;
        RECT  49.500 75.500 74.700 76.000 ;
        RECT  68.090 74.000 68.910 76.000 ;
        RECT  61.090 74.000 61.910 76.000 ;
        RECT  54.090 74.000 54.910 76.000 ;
        RECT  0.000 22.590 1.500 23.410 ;
        RECT  0.000 15.590 1.500 16.410 ;
        RECT  0.000 8.590 1.500 9.410 ;
        RECT  0.000 1.300 0.500 26.500 ;
        END
    END vdd
    PIN gnd
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M1 ;
        RECT  0.500 75.500 47.000 76.000 ;
        RECT  24.090 74.000 24.910 76.000 ;
        RECT  17.090 74.000 17.910 76.000 ;
        RECT  10.090 74.000 10.910 76.000 ;
        RECT  3.090 74.000 3.910 76.000 ;
        RECT  0.000 71.590 1.500 72.410 ;
        RECT  0.000 64.590 1.500 65.410 ;
        RECT  0.000 57.590 1.500 58.410 ;
        RECT  0.000 50.590 1.500 51.410 ;
        RECT  0.000 29.000 0.500 75.500 ;
        END
    END gnd
    OBS
        LAYER M1 ;
        RECT  2.090 1.300 31.000 7.000 ;
        RECT  2.090 11.000 31.000 14.000 ;
        RECT  2.090 18.000 31.000 21.000 ;
        RECT  2.090 25.000 31.000 49.000 ;
        RECT  2.090 53.000 31.000 56.000 ;
        RECT  2.090 60.000 31.000 63.000 ;
        RECT  2.090 67.000 31.000 70.000 ;
        RECT  3.090 1.300 31.000 72.410 ;
        RECT  32.500 2.800 73.200 72.410 ;
        RECT  5.500 1.300 8.500 73.910 ;
        RECT  12.500 1.300 15.500 73.910 ;
        RECT  19.500 1.300 22.500 73.910 ;
        RECT  26.500 1.300 31.000 73.910 ;
        RECT  32.500 2.800 52.500 73.910 ;
        RECT  56.500 2.800 59.500 73.910 ;
        RECT  63.500 2.800 66.500 73.910 ;
        RECT  70.500 2.800 73.200 73.910 ;
        RECT  73.200 43.525 73.250 73.910 ;
        RECT  73.250 43.575 73.300 73.910 ;
        RECT  73.300 43.625 73.350 73.910 ;
        RECT  73.350 43.675 73.400 73.910 ;
        RECT  73.400 43.725 73.450 73.910 ;
        RECT  73.450 43.775 73.500 73.910 ;
        RECT  73.500 43.825 73.550 73.910 ;
        RECT  73.550 43.875 73.600 73.910 ;
        RECT  73.600 43.925 73.650 73.910 ;
        RECT  73.650 43.975 73.700 73.910 ;
        RECT  73.700 44.025 73.750 73.910 ;
        RECT  73.750 44.075 73.800 73.910 ;
        RECT  73.800 44.125 73.850 73.910 ;
        RECT  73.850 44.175 73.900 73.910 ;
        RECT  73.900 44.225 73.950 73.910 ;
        RECT  73.950 44.275 74.000 73.910 ;
        RECT  74.000 44.325 74.050 73.910 ;
        RECT  74.050 44.375 74.100 73.910 ;
        RECT  74.100 44.425 74.150 73.910 ;
        RECT  74.150 44.475 74.200 73.910 ;
        RECT  74.200 44.525 74.250 73.910 ;
        RECT  74.250 44.575 74.300 73.910 ;
        RECT  74.300 44.625 74.350 73.910 ;
        RECT  74.350 44.675 74.400 73.910 ;
        RECT  74.400 44.725 74.450 73.910 ;
        RECT  74.450 44.775 74.500 73.910 ;
        RECT  74.500 44.825 74.550 73.910 ;
        RECT  74.550 44.875 74.600 73.910 ;
        RECT  74.600 44.925 74.650 73.910 ;
        RECT  74.650 44.975 74.700 73.910 ;
        RECT  31.000 1.325 31.050 73.910 ;
        RECT  31.050 1.375 31.100 73.910 ;
        RECT  31.100 1.425 31.150 73.910 ;
        RECT  31.150 1.475 31.200 73.910 ;
        RECT  31.200 1.525 31.250 73.910 ;
        RECT  31.250 1.575 31.300 73.910 ;
        RECT  31.300 1.625 31.350 73.910 ;
        RECT  31.350 1.675 31.400 73.910 ;
        RECT  31.400 1.725 31.450 73.910 ;
        RECT  31.450 1.775 31.500 73.910 ;
        RECT  31.500 1.825 31.550 73.910 ;
        RECT  31.550 1.875 31.600 73.910 ;
        RECT  31.600 1.925 31.650 73.910 ;
        RECT  31.650 1.975 31.700 73.910 ;
        RECT  31.700 2.025 31.750 73.910 ;
        RECT  31.750 2.075 31.800 73.910 ;
        RECT  31.800 2.125 31.850 73.910 ;
        RECT  31.850 2.175 31.900 73.910 ;
        RECT  31.900 2.225 31.950 73.910 ;
        RECT  31.950 2.275 32.000 73.910 ;
        RECT  32.000 2.325 32.050 73.910 ;
        RECT  32.050 2.375 32.100 73.910 ;
        RECT  32.100 2.425 32.150 73.910 ;
        RECT  32.150 2.475 32.200 73.910 ;
        RECT  32.200 2.525 32.250 73.910 ;
        RECT  32.250 2.575 32.300 73.910 ;
        RECT  32.300 2.625 32.350 73.910 ;
        RECT  32.350 2.675 32.400 73.910 ;
        RECT  32.400 2.725 32.450 73.910 ;
        RECT  32.450 2.775 32.500 73.910 ;
        LAYER M2 ;
        RECT  0.000 1.300 31.000 26.500 ;
        RECT  0.000 36.500 31.000 37.500 ;
        RECT  0.000 39.500 31.000 40.500 ;
        RECT  1.500 1.300 31.000 74.500 ;
        RECT  32.500 2.800 73.200 74.500 ;
        RECT  0.000 47.500 28.500 75.500 ;
        RECT  0.500 47.500 28.500 76.000 ;
        RECT  35.500 2.800 36.500 76.000 ;
        RECT  38.500 2.800 39.500 76.000 ;
        RECT  49.500 2.800 73.200 76.000 ;
        RECT  73.200 43.525 73.250 76.000 ;
        RECT  73.250 43.575 73.300 76.000 ;
        RECT  73.300 43.625 73.350 76.000 ;
        RECT  73.350 43.675 73.400 76.000 ;
        RECT  73.400 43.725 73.450 76.000 ;
        RECT  73.450 43.775 73.500 76.000 ;
        RECT  73.500 43.825 73.550 76.000 ;
        RECT  73.550 43.875 73.600 76.000 ;
        RECT  73.600 43.925 73.650 76.000 ;
        RECT  73.650 43.975 73.700 76.000 ;
        RECT  73.700 44.025 73.750 76.000 ;
        RECT  73.750 44.075 73.800 76.000 ;
        RECT  73.800 44.125 73.850 76.000 ;
        RECT  73.850 44.175 73.900 76.000 ;
        RECT  73.900 44.225 73.950 76.000 ;
        RECT  73.950 44.275 74.000 76.000 ;
        RECT  74.000 44.325 74.050 76.000 ;
        RECT  74.050 44.375 74.100 76.000 ;
        RECT  74.100 44.425 74.150 76.000 ;
        RECT  74.150 44.475 74.200 76.000 ;
        RECT  74.200 44.525 74.250 76.000 ;
        RECT  74.250 44.575 74.300 76.000 ;
        RECT  74.300 44.625 74.350 76.000 ;
        RECT  74.350 44.675 74.400 76.000 ;
        RECT  74.400 44.725 74.450 76.000 ;
        RECT  74.450 44.775 74.500 76.000 ;
        RECT  74.500 44.825 74.550 76.000 ;
        RECT  74.550 44.875 74.600 76.000 ;
        RECT  74.600 44.925 74.650 76.000 ;
        RECT  74.650 44.975 74.700 76.000 ;
        RECT  31.000 1.325 31.050 74.500 ;
        RECT  31.050 1.375 31.100 74.500 ;
        RECT  31.100 1.425 31.150 74.500 ;
        RECT  31.150 1.475 31.200 74.500 ;
        RECT  31.200 1.525 31.250 74.500 ;
        RECT  31.250 1.575 31.300 74.500 ;
        RECT  31.300 1.625 31.350 74.500 ;
        RECT  31.350 1.675 31.400 74.500 ;
        RECT  31.400 1.725 31.450 74.500 ;
        RECT  31.450 1.775 31.500 74.500 ;
        RECT  31.500 1.825 31.550 74.500 ;
        RECT  31.550 1.875 31.600 74.500 ;
        RECT  31.600 1.925 31.650 74.500 ;
        RECT  31.650 1.975 31.700 74.500 ;
        RECT  31.700 2.025 31.750 74.500 ;
        RECT  31.750 2.075 31.800 74.500 ;
        RECT  31.800 2.125 31.850 74.500 ;
        RECT  31.850 2.175 31.900 74.500 ;
        RECT  31.900 2.225 31.950 74.500 ;
        RECT  31.950 2.275 32.000 74.500 ;
        RECT  32.000 2.325 32.050 74.500 ;
        RECT  32.050 2.375 32.100 74.500 ;
        RECT  32.100 2.425 32.150 74.500 ;
        RECT  32.150 2.475 32.200 74.500 ;
        RECT  32.200 2.525 32.250 74.500 ;
        RECT  32.250 2.575 32.300 74.500 ;
        RECT  32.300 2.625 32.350 74.500 ;
        RECT  32.350 2.675 32.400 74.500 ;
        RECT  32.400 2.725 32.450 74.500 ;
        RECT  32.450 2.775 32.500 74.500 ;
        LAYER M3 ;
        RECT  1.500 2.800 73.200 74.500 ;
        LAYER M4 ;
        RECT  1.500 2.800 73.200 74.500 ;
        LAYER M5 ;
        RECT  1.500 2.800 73.200 74.500 ;
        LAYER M6 ;
        RECT  1.500 2.800 73.200 74.500 ;
        LAYER M7 ;
        RECT  1.500 2.800 73.200 74.500 ;
        LAYER AP ;
        RECT  1.000 2.300 73.700 75.000 ;
    END
END PADSPACE_C_74x74u_CH

MACRO PADSPACE_C_74x48u_CH_Rot
  CLASS ENDCAP BOTTOMLEFT ;
  ORIGIN 0 0 ;
  FOREIGN PADSPACE_C_74x48u_CH_Rot 0 0 ;
  SIZE 48 BY 76 ;
  SYMMETRY X Y R90 ;
  SITE IOSite ;
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 4.55 27.33 4.65 27.43 ;
        RECT 4.55 26.93 4.65 27.03 ;
        RECT 4.55 26.53 4.65 26.63 ;
        RECT 4.55 26.13 4.65 26.23 ;
        RECT 4.55 25.73 4.65 25.83 ;
        RECT 4.55 25.33 4.65 25.43 ;
        RECT 4.55 24.93 4.65 25.03 ;
        RECT 4.55 24.53 4.65 24.63 ;
        RECT 4.55 24.13 4.65 24.23 ;
        RECT 4.55 23.73 4.65 23.83 ;
        RECT 4.55 23.33 4.65 23.43 ;
        RECT 4.55 22.93 4.65 23.03 ;
        RECT 4.55 22.53 4.65 22.63 ;
        RECT 4.55 22.13 4.65 22.23 ;
        RECT 4.55 21.73 4.65 21.83 ;
        RECT 4.55 21.33 4.65 21.43 ;
        RECT 4.55 20.93 4.65 21.03 ;
        RECT 4.55 20.53 4.65 20.63 ;
        RECT 4.55 20.13 4.65 20.23 ;
        RECT 4.55 19.73 4.65 19.83 ;
        RECT 4.55 19.33 4.65 19.43 ;
        RECT 4.55 18.93 4.65 19.03 ;
        RECT 4.55 18.53 4.65 18.63 ;
        RECT 4.55 18.13 4.65 18.23 ;
        RECT 4.55 17.73 4.65 17.83 ;
        RECT 4.55 17.33 4.65 17.43 ;
        RECT 4.55 16.93 4.65 17.03 ;
        RECT 4.55 16.53 4.65 16.63 ;
        RECT 4.55 16.13 4.65 16.23 ;
        RECT 4.55 15.73 4.65 15.83 ;
        RECT 4.55 15.33 4.65 15.43 ;
        RECT 4.55 14.93 4.65 15.03 ;
        RECT 4.55 14.53 4.65 14.63 ;
        RECT 4.55 14.13 4.65 14.23 ;
        RECT 4.55 13.73 4.65 13.83 ;
        RECT 4.55 13.33 4.65 13.43 ;
        RECT 4.55 12.93 4.65 13.03 ;
        RECT 4.55 12.53 4.65 12.63 ;
        RECT 4.55 12.13 4.65 12.23 ;
        RECT 4.55 11.73 4.65 11.83 ;
        RECT 4.55 11.33 4.65 11.43 ;
        RECT 4.55 10.93 4.65 11.03 ;
        RECT 4.55 10.53 4.65 10.63 ;
        RECT 4.55 10.13 4.65 10.23 ;
        RECT 4.55 9.73 4.65 9.83 ;
        RECT 4.55 9.33 4.65 9.43 ;
        RECT 4.55 8.93 4.65 9.03 ;
        RECT 4.55 8.53 4.65 8.63 ;
        RECT 4.55 8.13 4.65 8.23 ;
        RECT 4.55 7.73 4.65 7.83 ;
        RECT 4.55 7.33 4.65 7.43 ;
        RECT 4.55 6.93 4.65 7.03 ;
        RECT 4.55 6.53 4.65 6.63 ;
        RECT 4.55 6.13 4.65 6.23 ;
        RECT 4.55 5.73 4.65 5.83 ;
        RECT 4.55 5.33 4.65 5.43 ;
        RECT 4.55 4.93 4.65 5.03 ;
        RECT 4.55 4.53 4.65 4.63 ;
        RECT 4.55 4.13 4.65 4.23 ;
        RECT 4.55 3.73 4.65 3.83 ;
        RECT 4.75 27.33 4.85 27.43 ;
        RECT 4.75 26.93 4.85 27.03 ;
        RECT 4.75 26.53 4.85 26.63 ;
        RECT 4.75 26.13 4.85 26.23 ;
        RECT 4.75 25.73 4.85 25.83 ;
        RECT 4.75 25.33 4.85 25.43 ;
        RECT 4.75 24.93 4.85 25.03 ;
        RECT 4.75 24.53 4.85 24.63 ;
        RECT 4.75 24.13 4.85 24.23 ;
        RECT 4.75 23.73 4.85 23.83 ;
        RECT 4.75 23.33 4.85 23.43 ;
        RECT 4.75 22.93 4.85 23.03 ;
        RECT 4.75 22.53 4.85 22.63 ;
        RECT 4.75 22.13 4.85 22.23 ;
        RECT 4.75 21.73 4.85 21.83 ;
        RECT 4.75 21.33 4.85 21.43 ;
        RECT 4.75 20.93 4.85 21.03 ;
        RECT 4.75 20.53 4.85 20.63 ;
        RECT 4.75 20.13 4.85 20.23 ;
        RECT 4.75 19.73 4.85 19.83 ;
        RECT 4.75 19.33 4.85 19.43 ;
        RECT 4.75 18.93 4.85 19.03 ;
        RECT 4.75 18.53 4.85 18.63 ;
        RECT 4.75 18.13 4.85 18.23 ;
        RECT 4.75 17.73 4.85 17.83 ;
        RECT 4.75 17.33 4.85 17.43 ;
        RECT 4.75 16.93 4.85 17.03 ;
        RECT 4.75 16.53 4.85 16.63 ;
        RECT 4.75 16.13 4.85 16.23 ;
        RECT 4.75 15.73 4.85 15.83 ;
        RECT 4.75 15.33 4.85 15.43 ;
        RECT 4.75 14.93 4.85 15.03 ;
        RECT 4.75 14.53 4.85 14.63 ;
        RECT 4.75 14.13 4.85 14.23 ;
        RECT 4.75 13.73 4.85 13.83 ;
        RECT 4.75 13.33 4.85 13.43 ;
        RECT 4.75 12.93 4.85 13.03 ;
        RECT 4.75 12.53 4.85 12.63 ;
        RECT 4.75 12.13 4.85 12.23 ;
        RECT 4.75 11.73 4.85 11.83 ;
        RECT 4.75 11.33 4.85 11.43 ;
        RECT 4.75 10.93 4.85 11.03 ;
        RECT 4.75 10.53 4.85 10.63 ;
        RECT 4.75 10.13 4.85 10.23 ;
        RECT 4.75 9.73 4.85 9.83 ;
        RECT 4.75 9.33 4.85 9.43 ;
        RECT 4.75 8.93 4.85 9.03 ;
        RECT 4.75 8.53 4.85 8.63 ;
        RECT 4.75 8.13 4.85 8.23 ;
        RECT 4.75 7.73 4.85 7.83 ;
        RECT 4.75 7.33 4.85 7.43 ;
        RECT 4.75 6.93 4.85 7.03 ;
        RECT 4.75 6.53 4.85 6.63 ;
        RECT 4.75 6.13 4.85 6.23 ;
        RECT 4.75 5.73 4.85 5.83 ;
        RECT 4.75 5.33 4.85 5.43 ;
        RECT 4.75 4.93 4.85 5.03 ;
        RECT 4.75 4.53 4.85 4.63 ;
        RECT 4.75 4.13 4.85 4.23 ;
        RECT 4.75 3.73 4.85 3.83 ;
        RECT 4.95 27.33 5.05 27.43 ;
        RECT 4.95 26.93 5.05 27.03 ;
        RECT 4.95 26.53 5.05 26.63 ;
        RECT 4.95 26.13 5.05 26.23 ;
        RECT 4.95 25.73 5.05 25.83 ;
        RECT 4.95 25.33 5.05 25.43 ;
        RECT 4.95 24.93 5.05 25.03 ;
        RECT 4.95 24.53 5.05 24.63 ;
        RECT 4.95 24.13 5.05 24.23 ;
        RECT 4.95 23.73 5.05 23.83 ;
        RECT 4.95 23.33 5.05 23.43 ;
        RECT 4.95 22.93 5.05 23.03 ;
        RECT 4.95 22.53 5.05 22.63 ;
        RECT 4.95 22.13 5.05 22.23 ;
        RECT 4.95 21.73 5.05 21.83 ;
        RECT 4.95 21.33 5.05 21.43 ;
        RECT 4.95 20.93 5.05 21.03 ;
        RECT 4.95 20.53 5.05 20.63 ;
        RECT 4.95 20.13 5.05 20.23 ;
        RECT 4.95 19.73 5.05 19.83 ;
        RECT 4.95 19.33 5.05 19.43 ;
        RECT 4.95 18.93 5.05 19.03 ;
        RECT 4.95 18.53 5.05 18.63 ;
        RECT 4.95 18.13 5.05 18.23 ;
        RECT 4.95 17.73 5.05 17.83 ;
        RECT 4.95 17.33 5.05 17.43 ;
        RECT 4.95 16.93 5.05 17.03 ;
        RECT 4.95 16.53 5.05 16.63 ;
        RECT 4.95 16.13 5.05 16.23 ;
        RECT 4.95 15.73 5.05 15.83 ;
        RECT 4.95 15.33 5.05 15.43 ;
        RECT 4.95 14.93 5.05 15.03 ;
        RECT 4.95 14.53 5.05 14.63 ;
        RECT 4.95 14.13 5.05 14.23 ;
        RECT 4.95 13.73 5.05 13.83 ;
        RECT 4.95 13.33 5.05 13.43 ;
        RECT 4.95 12.93 5.05 13.03 ;
        RECT 4.95 12.53 5.05 12.63 ;
        RECT 4.95 12.13 5.05 12.23 ;
        RECT 4.95 11.73 5.05 11.83 ;
        RECT 4.95 11.33 5.05 11.43 ;
        RECT 4.95 10.93 5.05 11.03 ;
        RECT 4.95 10.53 5.05 10.63 ;
        RECT 4.95 10.13 5.05 10.23 ;
        RECT 4.95 9.73 5.05 9.83 ;
        RECT 4.95 9.33 5.05 9.43 ;
        RECT 4.95 8.93 5.05 9.03 ;
        RECT 4.95 8.53 5.05 8.63 ;
        RECT 4.95 8.13 5.05 8.23 ;
        RECT 4.95 7.73 5.05 7.83 ;
        RECT 4.95 7.33 5.05 7.43 ;
        RECT 4.95 6.93 5.05 7.03 ;
        RECT 4.95 6.53 5.05 6.63 ;
        RECT 4.95 6.13 5.05 6.23 ;
        RECT 4.95 5.73 5.05 5.83 ;
        RECT 4.95 5.33 5.05 5.43 ;
        RECT 4.95 4.93 5.05 5.03 ;
        RECT 4.95 4.53 5.05 4.63 ;
        RECT 4.95 4.13 5.05 4.23 ;
        RECT 4.95 3.73 5.05 3.83 ;
        RECT 10.45 27.33 10.55 27.43 ;
        RECT 10.45 26.93 10.55 27.03 ;
        RECT 10.45 26.53 10.55 26.63 ;
        RECT 10.45 26.13 10.55 26.23 ;
        RECT 10.45 25.73 10.55 25.83 ;
        RECT 10.45 25.33 10.55 25.43 ;
        RECT 10.45 24.93 10.55 25.03 ;
        RECT 10.45 24.53 10.55 24.63 ;
        RECT 10.45 24.13 10.55 24.23 ;
        RECT 10.45 23.73 10.55 23.83 ;
        RECT 10.45 23.33 10.55 23.43 ;
        RECT 10.45 22.93 10.55 23.03 ;
        RECT 10.45 22.53 10.55 22.63 ;
        RECT 10.45 22.13 10.55 22.23 ;
        RECT 10.45 21.73 10.55 21.83 ;
        RECT 10.45 21.33 10.55 21.43 ;
        RECT 10.45 20.93 10.55 21.03 ;
        RECT 10.45 20.53 10.55 20.63 ;
        RECT 10.45 20.13 10.55 20.23 ;
        RECT 10.45 19.73 10.55 19.83 ;
        RECT 10.45 19.33 10.55 19.43 ;
        RECT 10.45 18.93 10.55 19.03 ;
        RECT 10.45 18.53 10.55 18.63 ;
        RECT 10.45 18.13 10.55 18.23 ;
        RECT 10.45 17.73 10.55 17.83 ;
        RECT 10.45 17.33 10.55 17.43 ;
        RECT 10.45 16.93 10.55 17.03 ;
        RECT 10.45 16.53 10.55 16.63 ;
        RECT 10.45 16.13 10.55 16.23 ;
        RECT 10.45 15.73 10.55 15.83 ;
        RECT 10.45 15.33 10.55 15.43 ;
        RECT 10.45 14.93 10.55 15.03 ;
        RECT 10.45 14.53 10.55 14.63 ;
        RECT 10.45 14.13 10.55 14.23 ;
        RECT 10.45 13.73 10.55 13.83 ;
        RECT 10.45 13.33 10.55 13.43 ;
        RECT 10.45 12.93 10.55 13.03 ;
        RECT 10.45 12.53 10.55 12.63 ;
        RECT 10.45 12.13 10.55 12.23 ;
        RECT 10.45 11.73 10.55 11.83 ;
        RECT 10.45 11.33 10.55 11.43 ;
        RECT 10.45 10.93 10.55 11.03 ;
        RECT 10.45 10.53 10.55 10.63 ;
        RECT 10.45 10.13 10.55 10.23 ;
        RECT 10.45 9.73 10.55 9.83 ;
        RECT 10.45 9.33 10.55 9.43 ;
        RECT 10.45 8.93 10.55 9.03 ;
        RECT 10.45 8.53 10.55 8.63 ;
        RECT 10.45 8.13 10.55 8.23 ;
        RECT 10.45 7.73 10.55 7.83 ;
        RECT 10.45 7.33 10.55 7.43 ;
        RECT 10.45 6.93 10.55 7.03 ;
        RECT 10.45 6.53 10.55 6.63 ;
        RECT 10.45 6.13 10.55 6.23 ;
        RECT 10.45 5.73 10.55 5.83 ;
        RECT 10.45 5.33 10.55 5.43 ;
        RECT 10.45 4.93 10.55 5.03 ;
        RECT 10.45 4.53 10.55 4.63 ;
        RECT 10.45 4.13 10.55 4.23 ;
        RECT 10.45 3.73 10.55 3.83 ;
        RECT 10.65 27.33 10.75 27.43 ;
        RECT 10.65 26.93 10.75 27.03 ;
        RECT 10.65 26.53 10.75 26.63 ;
        RECT 10.65 26.13 10.75 26.23 ;
        RECT 10.65 25.73 10.75 25.83 ;
        RECT 10.65 25.33 10.75 25.43 ;
        RECT 10.65 24.93 10.75 25.03 ;
        RECT 10.65 24.53 10.75 24.63 ;
        RECT 10.65 24.13 10.75 24.23 ;
        RECT 10.65 23.73 10.75 23.83 ;
        RECT 10.65 23.33 10.75 23.43 ;
        RECT 10.65 22.93 10.75 23.03 ;
        RECT 10.65 22.53 10.75 22.63 ;
        RECT 10.65 22.13 10.75 22.23 ;
        RECT 10.65 21.73 10.75 21.83 ;
        RECT 10.65 21.33 10.75 21.43 ;
        RECT 10.65 20.93 10.75 21.03 ;
        RECT 10.65 20.53 10.75 20.63 ;
        RECT 10.65 20.13 10.75 20.23 ;
        RECT 10.65 19.73 10.75 19.83 ;
        RECT 10.65 19.33 10.75 19.43 ;
        RECT 10.65 18.93 10.75 19.03 ;
        RECT 10.65 18.53 10.75 18.63 ;
        RECT 10.65 18.13 10.75 18.23 ;
        RECT 10.65 17.73 10.75 17.83 ;
        RECT 10.65 17.33 10.75 17.43 ;
        RECT 10.65 16.93 10.75 17.03 ;
        RECT 10.65 16.53 10.75 16.63 ;
        RECT 10.65 16.13 10.75 16.23 ;
        RECT 10.65 15.73 10.75 15.83 ;
        RECT 10.65 15.33 10.75 15.43 ;
        RECT 10.65 14.93 10.75 15.03 ;
        RECT 10.65 14.53 10.75 14.63 ;
        RECT 10.65 14.13 10.75 14.23 ;
        RECT 10.65 13.73 10.75 13.83 ;
        RECT 10.65 13.33 10.75 13.43 ;
        RECT 10.65 12.93 10.75 13.03 ;
        RECT 10.65 12.53 10.75 12.63 ;
        RECT 10.65 12.13 10.75 12.23 ;
        RECT 10.65 11.73 10.75 11.83 ;
        RECT 10.65 11.33 10.75 11.43 ;
        RECT 10.65 10.93 10.75 11.03 ;
        RECT 10.65 10.53 10.75 10.63 ;
        RECT 10.65 10.13 10.75 10.23 ;
        RECT 10.65 9.73 10.75 9.83 ;
        RECT 10.65 9.33 10.75 9.43 ;
        RECT 10.65 8.93 10.75 9.03 ;
        RECT 10.65 8.53 10.75 8.63 ;
        RECT 10.65 8.13 10.75 8.23 ;
        RECT 10.65 7.73 10.75 7.83 ;
        RECT 10.65 7.33 10.75 7.43 ;
        RECT 10.65 6.93 10.75 7.03 ;
        RECT 10.65 6.53 10.75 6.63 ;
        RECT 10.65 6.13 10.75 6.23 ;
        RECT 10.65 5.73 10.75 5.83 ;
        RECT 10.65 5.33 10.75 5.43 ;
        RECT 10.65 4.93 10.75 5.03 ;
        RECT 10.65 4.53 10.75 4.63 ;
        RECT 10.65 4.13 10.75 4.23 ;
        RECT 10.65 3.73 10.75 3.83 ;
        RECT 10.85 27.33 10.95 27.43 ;
        RECT 10.85 26.93 10.95 27.03 ;
        RECT 10.85 26.53 10.95 26.63 ;
        RECT 10.85 26.13 10.95 26.23 ;
        RECT 10.85 25.73 10.95 25.83 ;
        RECT 10.85 25.33 10.95 25.43 ;
        RECT 10.85 24.93 10.95 25.03 ;
        RECT 10.85 24.53 10.95 24.63 ;
        RECT 10.85 24.13 10.95 24.23 ;
        RECT 10.85 23.73 10.95 23.83 ;
        RECT 10.85 23.33 10.95 23.43 ;
        RECT 10.85 22.93 10.95 23.03 ;
        RECT 10.85 22.53 10.95 22.63 ;
        RECT 10.85 22.13 10.95 22.23 ;
        RECT 10.85 21.73 10.95 21.83 ;
        RECT 10.85 21.33 10.95 21.43 ;
        RECT 10.85 20.93 10.95 21.03 ;
        RECT 10.85 20.53 10.95 20.63 ;
        RECT 10.85 20.13 10.95 20.23 ;
        RECT 10.85 19.73 10.95 19.83 ;
        RECT 10.85 19.33 10.95 19.43 ;
        RECT 10.85 18.93 10.95 19.03 ;
        RECT 10.85 18.53 10.95 18.63 ;
        RECT 10.85 18.13 10.95 18.23 ;
        RECT 10.85 17.73 10.95 17.83 ;
        RECT 10.85 17.33 10.95 17.43 ;
        RECT 10.85 16.93 10.95 17.03 ;
        RECT 10.85 16.53 10.95 16.63 ;
        RECT 10.85 16.13 10.95 16.23 ;
        RECT 10.85 15.73 10.95 15.83 ;
        RECT 10.85 15.33 10.95 15.43 ;
        RECT 10.85 14.93 10.95 15.03 ;
        RECT 10.85 14.53 10.95 14.63 ;
        RECT 10.85 14.13 10.95 14.23 ;
        RECT 10.85 13.73 10.95 13.83 ;
        RECT 10.85 13.33 10.95 13.43 ;
        RECT 10.85 12.93 10.95 13.03 ;
        RECT 10.85 12.53 10.95 12.63 ;
        RECT 10.85 12.13 10.95 12.23 ;
        RECT 10.85 11.73 10.95 11.83 ;
        RECT 10.85 11.33 10.95 11.43 ;
        RECT 10.85 10.93 10.95 11.03 ;
        RECT 10.85 10.53 10.95 10.63 ;
        RECT 10.85 10.13 10.95 10.23 ;
        RECT 10.85 9.73 10.95 9.83 ;
        RECT 10.85 9.33 10.95 9.43 ;
        RECT 10.85 8.93 10.95 9.03 ;
        RECT 10.85 8.53 10.95 8.63 ;
        RECT 10.85 8.13 10.95 8.23 ;
        RECT 10.85 7.73 10.95 7.83 ;
        RECT 10.85 7.33 10.95 7.43 ;
        RECT 10.85 6.93 10.95 7.03 ;
        RECT 10.85 6.53 10.95 6.63 ;
        RECT 10.85 6.13 10.95 6.23 ;
        RECT 10.85 5.73 10.95 5.83 ;
        RECT 10.85 5.33 10.95 5.43 ;
        RECT 10.85 4.93 10.95 5.03 ;
        RECT 10.85 4.53 10.95 4.63 ;
        RECT 10.85 4.13 10.95 4.23 ;
        RECT 10.85 3.73 10.95 3.83 ;
        RECT 11.05 27.33 11.15 27.43 ;
        RECT 11.05 26.93 11.15 27.03 ;
        RECT 11.05 26.53 11.15 26.63 ;
        RECT 11.05 26.13 11.15 26.23 ;
        RECT 11.05 25.73 11.15 25.83 ;
        RECT 11.05 25.33 11.15 25.43 ;
        RECT 11.05 24.93 11.15 25.03 ;
        RECT 11.05 24.53 11.15 24.63 ;
        RECT 11.05 24.13 11.15 24.23 ;
        RECT 11.05 23.73 11.15 23.83 ;
        RECT 11.05 23.33 11.15 23.43 ;
        RECT 11.05 22.93 11.15 23.03 ;
        RECT 11.05 22.53 11.15 22.63 ;
        RECT 11.05 22.13 11.15 22.23 ;
        RECT 11.05 21.73 11.15 21.83 ;
        RECT 11.05 21.33 11.15 21.43 ;
        RECT 11.05 20.93 11.15 21.03 ;
        RECT 11.05 20.53 11.15 20.63 ;
        RECT 11.05 20.13 11.15 20.23 ;
        RECT 11.05 19.73 11.15 19.83 ;
        RECT 11.05 19.33 11.15 19.43 ;
        RECT 11.05 18.93 11.15 19.03 ;
        RECT 11.05 18.53 11.15 18.63 ;
        RECT 11.05 18.13 11.15 18.23 ;
        RECT 11.05 17.73 11.15 17.83 ;
        RECT 11.05 17.33 11.15 17.43 ;
        RECT 11.05 16.93 11.15 17.03 ;
        RECT 11.05 16.53 11.15 16.63 ;
        RECT 11.05 16.13 11.15 16.23 ;
        RECT 11.05 15.73 11.15 15.83 ;
        RECT 11.05 15.33 11.15 15.43 ;
        RECT 11.05 14.93 11.15 15.03 ;
        RECT 11.05 14.53 11.15 14.63 ;
        RECT 11.05 14.13 11.15 14.23 ;
        RECT 11.05 13.73 11.15 13.83 ;
        RECT 11.05 13.33 11.15 13.43 ;
        RECT 11.05 12.93 11.15 13.03 ;
        RECT 11.05 12.53 11.15 12.63 ;
        RECT 11.05 12.13 11.15 12.23 ;
        RECT 11.05 11.73 11.15 11.83 ;
        RECT 11.05 11.33 11.15 11.43 ;
        RECT 11.05 10.93 11.15 11.03 ;
        RECT 11.05 10.53 11.15 10.63 ;
        RECT 11.05 10.13 11.15 10.23 ;
        RECT 11.05 9.73 11.15 9.83 ;
        RECT 11.05 9.33 11.15 9.43 ;
        RECT 11.05 8.93 11.15 9.03 ;
        RECT 11.05 8.53 11.15 8.63 ;
        RECT 11.05 8.13 11.15 8.23 ;
        RECT 11.05 7.73 11.15 7.83 ;
        RECT 11.05 7.33 11.15 7.43 ;
        RECT 11.05 6.93 11.15 7.03 ;
        RECT 11.05 6.53 11.15 6.63 ;
        RECT 11.05 6.13 11.15 6.23 ;
        RECT 11.05 5.73 11.15 5.83 ;
        RECT 11.05 5.33 11.15 5.43 ;
        RECT 11.05 4.93 11.15 5.03 ;
        RECT 11.05 4.53 11.15 4.63 ;
        RECT 11.05 4.13 11.15 4.23 ;
        RECT 11.05 3.73 11.15 3.83 ;
        RECT 11.25 27.33 11.35 27.43 ;
        RECT 11.25 26.93 11.35 27.03 ;
        RECT 11.25 26.53 11.35 26.63 ;
        RECT 11.25 26.13 11.35 26.23 ;
        RECT 11.25 25.73 11.35 25.83 ;
        RECT 11.25 25.33 11.35 25.43 ;
        RECT 11.25 24.93 11.35 25.03 ;
        RECT 11.25 24.53 11.35 24.63 ;
        RECT 11.25 24.13 11.35 24.23 ;
        RECT 11.25 23.73 11.35 23.83 ;
        RECT 11.25 23.33 11.35 23.43 ;
        RECT 11.25 22.93 11.35 23.03 ;
        RECT 11.25 22.53 11.35 22.63 ;
        RECT 11.25 22.13 11.35 22.23 ;
        RECT 11.25 21.73 11.35 21.83 ;
        RECT 11.25 21.33 11.35 21.43 ;
        RECT 11.25 20.93 11.35 21.03 ;
        RECT 11.25 20.53 11.35 20.63 ;
        RECT 11.25 20.13 11.35 20.23 ;
        RECT 11.25 19.73 11.35 19.83 ;
        RECT 11.25 19.33 11.35 19.43 ;
        RECT 11.25 18.93 11.35 19.03 ;
        RECT 11.25 18.53 11.35 18.63 ;
        RECT 11.25 18.13 11.35 18.23 ;
        RECT 11.25 17.73 11.35 17.83 ;
        RECT 11.25 17.33 11.35 17.43 ;
        RECT 11.25 16.93 11.35 17.03 ;
        RECT 11.25 16.53 11.35 16.63 ;
        RECT 11.25 16.13 11.35 16.23 ;
        RECT 11.25 15.73 11.35 15.83 ;
        RECT 11.25 15.33 11.35 15.43 ;
        RECT 11.25 14.93 11.35 15.03 ;
        RECT 11.25 14.53 11.35 14.63 ;
        RECT 11.25 14.13 11.35 14.23 ;
        RECT 11.25 13.73 11.35 13.83 ;
        RECT 11.25 13.33 11.35 13.43 ;
        RECT 11.25 12.93 11.35 13.03 ;
        RECT 11.25 12.53 11.35 12.63 ;
        RECT 11.25 12.13 11.35 12.23 ;
        RECT 11.25 11.73 11.35 11.83 ;
        RECT 11.25 11.33 11.35 11.43 ;
        RECT 11.25 10.93 11.35 11.03 ;
        RECT 11.25 10.53 11.35 10.63 ;
        RECT 11.25 10.13 11.35 10.23 ;
        RECT 11.25 9.73 11.35 9.83 ;
        RECT 11.25 9.33 11.35 9.43 ;
        RECT 11.25 8.93 11.35 9.03 ;
        RECT 11.25 8.53 11.35 8.63 ;
        RECT 11.25 8.13 11.35 8.23 ;
        RECT 11.25 7.73 11.35 7.83 ;
        RECT 11.25 7.33 11.35 7.43 ;
        RECT 11.25 6.93 11.35 7.03 ;
        RECT 11.25 6.53 11.35 6.63 ;
        RECT 11.25 6.13 11.35 6.23 ;
        RECT 11.25 5.73 11.35 5.83 ;
        RECT 11.25 5.33 11.35 5.43 ;
        RECT 11.25 4.93 11.35 5.03 ;
        RECT 11.25 4.53 11.35 4.63 ;
        RECT 11.25 4.13 11.35 4.23 ;
        RECT 11.25 3.73 11.35 3.83 ;
        RECT 11.45 27.33 11.55 27.43 ;
        RECT 11.45 26.93 11.55 27.03 ;
        RECT 11.45 26.53 11.55 26.63 ;
        RECT 11.45 26.13 11.55 26.23 ;
        RECT 11.45 25.73 11.55 25.83 ;
        RECT 11.45 25.33 11.55 25.43 ;
        RECT 11.45 24.93 11.55 25.03 ;
        RECT 11.45 24.53 11.55 24.63 ;
        RECT 11.45 24.13 11.55 24.23 ;
        RECT 11.45 23.73 11.55 23.83 ;
        RECT 11.45 23.33 11.55 23.43 ;
        RECT 11.45 22.93 11.55 23.03 ;
        RECT 11.45 22.53 11.55 22.63 ;
        RECT 11.45 22.13 11.55 22.23 ;
        RECT 11.45 21.73 11.55 21.83 ;
        RECT 11.45 21.33 11.55 21.43 ;
        RECT 11.45 20.93 11.55 21.03 ;
        RECT 11.45 20.53 11.55 20.63 ;
        RECT 11.45 20.13 11.55 20.23 ;
        RECT 11.45 19.73 11.55 19.83 ;
        RECT 11.45 19.33 11.55 19.43 ;
        RECT 11.45 18.93 11.55 19.03 ;
        RECT 11.45 18.53 11.55 18.63 ;
        RECT 11.45 18.13 11.55 18.23 ;
        RECT 11.45 17.73 11.55 17.83 ;
        RECT 11.45 17.33 11.55 17.43 ;
        RECT 11.45 16.93 11.55 17.03 ;
        RECT 11.45 16.53 11.55 16.63 ;
        RECT 11.45 16.13 11.55 16.23 ;
        RECT 11.45 15.73 11.55 15.83 ;
        RECT 11.45 15.33 11.55 15.43 ;
        RECT 11.45 14.93 11.55 15.03 ;
        RECT 11.45 14.53 11.55 14.63 ;
        RECT 11.45 14.13 11.55 14.23 ;
        RECT 11.45 13.73 11.55 13.83 ;
        RECT 11.45 13.33 11.55 13.43 ;
        RECT 11.45 12.93 11.55 13.03 ;
        RECT 11.45 12.53 11.55 12.63 ;
        RECT 11.45 12.13 11.55 12.23 ;
        RECT 11.45 11.73 11.55 11.83 ;
        RECT 11.45 11.33 11.55 11.43 ;
        RECT 11.45 10.93 11.55 11.03 ;
        RECT 11.45 10.53 11.55 10.63 ;
        RECT 11.45 10.13 11.55 10.23 ;
        RECT 11.45 9.73 11.55 9.83 ;
        RECT 11.45 9.33 11.55 9.43 ;
        RECT 11.45 8.93 11.55 9.03 ;
        RECT 11.45 8.53 11.55 8.63 ;
        RECT 11.45 8.13 11.55 8.23 ;
        RECT 11.45 7.73 11.55 7.83 ;
        RECT 11.45 7.33 11.55 7.43 ;
        RECT 11.45 6.93 11.55 7.03 ;
        RECT 11.45 6.53 11.55 6.63 ;
        RECT 11.45 6.13 11.55 6.23 ;
        RECT 11.45 5.73 11.55 5.83 ;
        RECT 11.45 5.33 11.55 5.43 ;
        RECT 11.45 4.93 11.55 5.03 ;
        RECT 11.45 4.53 11.55 4.63 ;
        RECT 11.45 4.13 11.55 4.23 ;
        RECT 11.45 3.73 11.55 3.83 ;
        RECT 17.45 27.33 17.55 27.43 ;
        RECT 17.45 26.93 17.55 27.03 ;
        RECT 17.45 26.53 17.55 26.63 ;
        RECT 17.45 26.13 17.55 26.23 ;
        RECT 17.45 25.73 17.55 25.83 ;
        RECT 17.45 25.33 17.55 25.43 ;
        RECT 17.45 24.93 17.55 25.03 ;
        RECT 17.45 24.53 17.55 24.63 ;
        RECT 17.45 24.13 17.55 24.23 ;
        RECT 17.45 23.73 17.55 23.83 ;
        RECT 17.45 23.33 17.55 23.43 ;
        RECT 17.45 22.93 17.55 23.03 ;
        RECT 17.45 22.53 17.55 22.63 ;
        RECT 17.45 22.13 17.55 22.23 ;
        RECT 17.45 21.73 17.55 21.83 ;
        RECT 17.45 21.33 17.55 21.43 ;
        RECT 17.45 20.93 17.55 21.03 ;
        RECT 17.45 20.53 17.55 20.63 ;
        RECT 17.45 20.13 17.55 20.23 ;
        RECT 17.45 19.73 17.55 19.83 ;
        RECT 17.45 19.33 17.55 19.43 ;
        RECT 17.45 18.93 17.55 19.03 ;
        RECT 17.45 18.53 17.55 18.63 ;
        RECT 17.45 18.13 17.55 18.23 ;
        RECT 17.45 17.73 17.55 17.83 ;
        RECT 17.45 17.33 17.55 17.43 ;
        RECT 17.45 16.93 17.55 17.03 ;
        RECT 17.45 16.53 17.55 16.63 ;
        RECT 17.45 16.13 17.55 16.23 ;
        RECT 17.45 15.73 17.55 15.83 ;
        RECT 17.45 15.33 17.55 15.43 ;
        RECT 17.45 14.93 17.55 15.03 ;
        RECT 17.45 14.53 17.55 14.63 ;
        RECT 17.45 14.13 17.55 14.23 ;
        RECT 17.45 13.73 17.55 13.83 ;
        RECT 17.45 13.33 17.55 13.43 ;
        RECT 17.45 12.93 17.55 13.03 ;
        RECT 17.45 12.53 17.55 12.63 ;
        RECT 17.45 12.13 17.55 12.23 ;
        RECT 17.45 11.73 17.55 11.83 ;
        RECT 17.45 11.33 17.55 11.43 ;
        RECT 17.45 10.93 17.55 11.03 ;
        RECT 17.45 10.53 17.55 10.63 ;
        RECT 17.45 10.13 17.55 10.23 ;
        RECT 17.45 9.73 17.55 9.83 ;
        RECT 17.45 9.33 17.55 9.43 ;
        RECT 17.45 8.93 17.55 9.03 ;
        RECT 17.45 8.53 17.55 8.63 ;
        RECT 17.45 8.13 17.55 8.23 ;
        RECT 17.45 7.73 17.55 7.83 ;
        RECT 17.45 7.33 17.55 7.43 ;
        RECT 17.45 6.93 17.55 7.03 ;
        RECT 17.45 6.53 17.55 6.63 ;
        RECT 17.45 6.13 17.55 6.23 ;
        RECT 17.45 5.73 17.55 5.83 ;
        RECT 17.45 5.33 17.55 5.43 ;
        RECT 17.45 4.93 17.55 5.03 ;
        RECT 17.45 4.53 17.55 4.63 ;
        RECT 17.45 4.13 17.55 4.23 ;
        RECT 17.45 3.73 17.55 3.83 ;
        RECT 17.65 27.33 17.75 27.43 ;
        RECT 17.65 26.93 17.75 27.03 ;
        RECT 17.65 26.53 17.75 26.63 ;
        RECT 17.65 26.13 17.75 26.23 ;
        RECT 17.65 25.73 17.75 25.83 ;
        RECT 17.65 25.33 17.75 25.43 ;
        RECT 17.65 24.93 17.75 25.03 ;
        RECT 17.65 24.53 17.75 24.63 ;
        RECT 17.65 24.13 17.75 24.23 ;
        RECT 17.65 23.73 17.75 23.83 ;
        RECT 17.65 23.33 17.75 23.43 ;
        RECT 17.65 22.93 17.75 23.03 ;
        RECT 17.65 22.53 17.75 22.63 ;
        RECT 17.65 22.13 17.75 22.23 ;
        RECT 17.65 21.73 17.75 21.83 ;
        RECT 17.65 21.33 17.75 21.43 ;
        RECT 17.65 20.93 17.75 21.03 ;
        RECT 17.65 20.53 17.75 20.63 ;
        RECT 17.65 20.13 17.75 20.23 ;
        RECT 17.65 19.73 17.75 19.83 ;
        RECT 17.65 19.33 17.75 19.43 ;
        RECT 17.65 18.93 17.75 19.03 ;
        RECT 17.65 18.53 17.75 18.63 ;
        RECT 17.65 18.13 17.75 18.23 ;
        RECT 17.65 17.73 17.75 17.83 ;
        RECT 17.65 17.33 17.75 17.43 ;
        RECT 17.65 16.93 17.75 17.03 ;
        RECT 17.65 16.53 17.75 16.63 ;
        RECT 17.65 16.13 17.75 16.23 ;
        RECT 17.65 15.73 17.75 15.83 ;
        RECT 17.65 15.33 17.75 15.43 ;
        RECT 17.65 14.93 17.75 15.03 ;
        RECT 17.65 14.53 17.75 14.63 ;
        RECT 17.65 14.13 17.75 14.23 ;
        RECT 17.65 13.73 17.75 13.83 ;
        RECT 17.65 13.33 17.75 13.43 ;
        RECT 17.65 12.93 17.75 13.03 ;
        RECT 17.65 12.53 17.75 12.63 ;
        RECT 17.65 12.13 17.75 12.23 ;
        RECT 17.65 11.73 17.75 11.83 ;
        RECT 17.65 11.33 17.75 11.43 ;
        RECT 17.65 10.93 17.75 11.03 ;
        RECT 17.65 10.53 17.75 10.63 ;
        RECT 17.65 10.13 17.75 10.23 ;
        RECT 17.65 9.73 17.75 9.83 ;
        RECT 17.65 9.33 17.75 9.43 ;
        RECT 17.65 8.93 17.75 9.03 ;
        RECT 17.65 8.53 17.75 8.63 ;
        RECT 17.65 8.13 17.75 8.23 ;
        RECT 17.65 7.73 17.75 7.83 ;
        RECT 17.65 7.33 17.75 7.43 ;
        RECT 17.65 6.93 17.75 7.03 ;
        RECT 17.65 6.53 17.75 6.63 ;
        RECT 17.65 6.13 17.75 6.23 ;
        RECT 17.65 5.73 17.75 5.83 ;
        RECT 17.65 5.33 17.75 5.43 ;
        RECT 17.65 4.93 17.75 5.03 ;
        RECT 17.65 4.53 17.75 4.63 ;
        RECT 17.65 4.13 17.75 4.23 ;
        RECT 17.65 3.73 17.75 3.83 ;
        RECT 17.85 27.33 17.95 27.43 ;
        RECT 17.85 26.93 17.95 27.03 ;
        RECT 17.85 26.53 17.95 26.63 ;
        RECT 17.85 26.13 17.95 26.23 ;
        RECT 17.85 25.73 17.95 25.83 ;
        RECT 17.85 25.33 17.95 25.43 ;
        RECT 17.85 24.93 17.95 25.03 ;
        RECT 17.85 24.53 17.95 24.63 ;
        RECT 17.85 24.13 17.95 24.23 ;
        RECT 17.85 23.73 17.95 23.83 ;
        RECT 17.85 23.33 17.95 23.43 ;
        RECT 17.85 22.93 17.95 23.03 ;
        RECT 17.85 22.53 17.95 22.63 ;
        RECT 17.85 22.13 17.95 22.23 ;
        RECT 17.85 21.73 17.95 21.83 ;
        RECT 17.85 21.33 17.95 21.43 ;
        RECT 17.85 20.93 17.95 21.03 ;
        RECT 17.85 20.53 17.95 20.63 ;
        RECT 17.85 20.13 17.95 20.23 ;
        RECT 17.85 19.73 17.95 19.83 ;
        RECT 17.85 19.33 17.95 19.43 ;
        RECT 17.85 18.93 17.95 19.03 ;
        RECT 17.85 18.53 17.95 18.63 ;
        RECT 17.85 18.13 17.95 18.23 ;
        RECT 17.85 17.73 17.95 17.83 ;
        RECT 17.85 17.33 17.95 17.43 ;
        RECT 17.85 16.93 17.95 17.03 ;
        RECT 17.85 16.53 17.95 16.63 ;
        RECT 17.85 16.13 17.95 16.23 ;
        RECT 17.85 15.73 17.95 15.83 ;
        RECT 17.85 15.33 17.95 15.43 ;
        RECT 17.85 14.93 17.95 15.03 ;
        RECT 17.85 14.53 17.95 14.63 ;
        RECT 17.85 14.13 17.95 14.23 ;
        RECT 17.85 13.73 17.95 13.83 ;
        RECT 17.85 13.33 17.95 13.43 ;
        RECT 17.85 12.93 17.95 13.03 ;
        RECT 17.85 12.53 17.95 12.63 ;
        RECT 17.85 12.13 17.95 12.23 ;
        RECT 17.85 11.73 17.95 11.83 ;
        RECT 17.85 11.33 17.95 11.43 ;
        RECT 17.85 10.93 17.95 11.03 ;
        RECT 17.85 10.53 17.95 10.63 ;
        RECT 17.85 10.13 17.95 10.23 ;
        RECT 17.85 9.73 17.95 9.83 ;
        RECT 17.85 9.33 17.95 9.43 ;
        RECT 17.85 8.93 17.95 9.03 ;
        RECT 17.85 8.53 17.95 8.63 ;
        RECT 17.85 8.13 17.95 8.23 ;
        RECT 17.85 7.73 17.95 7.83 ;
        RECT 17.85 7.33 17.95 7.43 ;
        RECT 17.85 6.93 17.95 7.03 ;
        RECT 17.85 6.53 17.95 6.63 ;
        RECT 17.85 6.13 17.95 6.23 ;
        RECT 17.85 5.73 17.95 5.83 ;
        RECT 17.85 5.33 17.95 5.43 ;
        RECT 17.85 4.93 17.95 5.03 ;
        RECT 17.85 4.53 17.95 4.63 ;
        RECT 17.85 4.13 17.95 4.23 ;
        RECT 17.85 3.73 17.95 3.83 ;
        RECT 18.05 27.33 18.15 27.43 ;
        RECT 18.05 26.93 18.15 27.03 ;
        RECT 18.05 26.53 18.15 26.63 ;
        RECT 18.05 26.13 18.15 26.23 ;
        RECT 18.05 25.73 18.15 25.83 ;
        RECT 18.05 25.33 18.15 25.43 ;
        RECT 18.05 24.93 18.15 25.03 ;
        RECT 18.05 24.53 18.15 24.63 ;
        RECT 18.05 24.13 18.15 24.23 ;
        RECT 18.05 23.73 18.15 23.83 ;
        RECT 18.05 23.33 18.15 23.43 ;
        RECT 18.05 22.93 18.15 23.03 ;
        RECT 18.05 22.53 18.15 22.63 ;
        RECT 18.05 22.13 18.15 22.23 ;
        RECT 18.05 21.73 18.15 21.83 ;
        RECT 18.05 21.33 18.15 21.43 ;
        RECT 18.05 20.93 18.15 21.03 ;
        RECT 18.05 20.53 18.15 20.63 ;
        RECT 18.05 20.13 18.15 20.23 ;
        RECT 18.05 19.73 18.15 19.83 ;
        RECT 18.05 19.33 18.15 19.43 ;
        RECT 18.05 18.93 18.15 19.03 ;
        RECT 18.05 18.53 18.15 18.63 ;
        RECT 18.05 18.13 18.15 18.23 ;
        RECT 18.05 17.73 18.15 17.83 ;
        RECT 18.05 17.33 18.15 17.43 ;
        RECT 18.05 16.93 18.15 17.03 ;
        RECT 18.05 16.53 18.15 16.63 ;
        RECT 18.05 16.13 18.15 16.23 ;
        RECT 18.05 15.73 18.15 15.83 ;
        RECT 18.05 15.33 18.15 15.43 ;
        RECT 18.05 14.93 18.15 15.03 ;
        RECT 18.05 14.53 18.15 14.63 ;
        RECT 18.05 14.13 18.15 14.23 ;
        RECT 18.05 13.73 18.15 13.83 ;
        RECT 18.05 13.33 18.15 13.43 ;
        RECT 18.05 12.93 18.15 13.03 ;
        RECT 18.05 12.53 18.15 12.63 ;
        RECT 18.05 12.13 18.15 12.23 ;
        RECT 18.05 11.73 18.15 11.83 ;
        RECT 18.05 11.33 18.15 11.43 ;
        RECT 18.05 10.93 18.15 11.03 ;
        RECT 18.05 10.53 18.15 10.63 ;
        RECT 18.05 10.13 18.15 10.23 ;
        RECT 18.05 9.73 18.15 9.83 ;
        RECT 18.05 9.33 18.15 9.43 ;
        RECT 18.05 8.93 18.15 9.03 ;
        RECT 18.05 8.53 18.15 8.63 ;
        RECT 18.05 8.13 18.15 8.23 ;
        RECT 18.05 7.73 18.15 7.83 ;
        RECT 18.05 7.33 18.15 7.43 ;
        RECT 18.05 6.93 18.15 7.03 ;
        RECT 18.05 6.53 18.15 6.63 ;
        RECT 18.05 6.13 18.15 6.23 ;
        RECT 18.05 5.73 18.15 5.83 ;
        RECT 18.05 5.33 18.15 5.43 ;
        RECT 18.05 4.93 18.15 5.03 ;
        RECT 18.05 4.53 18.15 4.63 ;
        RECT 18.05 4.13 18.15 4.23 ;
        RECT 18.05 3.73 18.15 3.83 ;
        RECT 18.25 27.33 18.35 27.43 ;
        RECT 18.25 26.93 18.35 27.03 ;
        RECT 18.25 26.53 18.35 26.63 ;
        RECT 18.25 26.13 18.35 26.23 ;
        RECT 18.25 25.73 18.35 25.83 ;
        RECT 18.25 25.33 18.35 25.43 ;
        RECT 18.25 24.93 18.35 25.03 ;
        RECT 18.25 24.53 18.35 24.63 ;
        RECT 18.25 24.13 18.35 24.23 ;
        RECT 18.25 23.73 18.35 23.83 ;
        RECT 18.25 23.33 18.35 23.43 ;
        RECT 18.25 22.93 18.35 23.03 ;
        RECT 18.25 22.53 18.35 22.63 ;
        RECT 18.25 22.13 18.35 22.23 ;
        RECT 18.25 21.73 18.35 21.83 ;
        RECT 18.25 21.33 18.35 21.43 ;
        RECT 18.25 20.93 18.35 21.03 ;
        RECT 18.25 20.53 18.35 20.63 ;
        RECT 18.25 20.13 18.35 20.23 ;
        RECT 18.25 19.73 18.35 19.83 ;
        RECT 18.25 19.33 18.35 19.43 ;
        RECT 18.25 18.93 18.35 19.03 ;
        RECT 18.25 18.53 18.35 18.63 ;
        RECT 18.25 18.13 18.35 18.23 ;
        RECT 18.25 17.73 18.35 17.83 ;
        RECT 18.25 17.33 18.35 17.43 ;
        RECT 18.25 16.93 18.35 17.03 ;
        RECT 18.25 16.53 18.35 16.63 ;
        RECT 18.25 16.13 18.35 16.23 ;
        RECT 18.25 15.73 18.35 15.83 ;
        RECT 18.25 15.33 18.35 15.43 ;
        RECT 18.25 14.93 18.35 15.03 ;
        RECT 18.25 14.53 18.35 14.63 ;
        RECT 18.25 14.13 18.35 14.23 ;
        RECT 18.25 13.73 18.35 13.83 ;
        RECT 18.25 13.33 18.35 13.43 ;
        RECT 18.25 12.93 18.35 13.03 ;
        RECT 18.25 12.53 18.35 12.63 ;
        RECT 18.25 12.13 18.35 12.23 ;
        RECT 18.25 11.73 18.35 11.83 ;
        RECT 18.25 11.33 18.35 11.43 ;
        RECT 18.25 10.93 18.35 11.03 ;
        RECT 18.25 10.53 18.35 10.63 ;
        RECT 18.25 10.13 18.35 10.23 ;
        RECT 18.25 9.73 18.35 9.83 ;
        RECT 18.25 9.33 18.35 9.43 ;
        RECT 18.25 8.93 18.35 9.03 ;
        RECT 18.25 8.53 18.35 8.63 ;
        RECT 18.25 8.13 18.35 8.23 ;
        RECT 18.25 7.73 18.35 7.83 ;
        RECT 18.25 7.33 18.35 7.43 ;
        RECT 18.25 6.93 18.35 7.03 ;
        RECT 18.25 6.53 18.35 6.63 ;
        RECT 18.25 6.13 18.35 6.23 ;
        RECT 18.25 5.73 18.35 5.83 ;
        RECT 18.25 5.33 18.35 5.43 ;
        RECT 18.25 4.93 18.35 5.03 ;
        RECT 18.25 4.53 18.35 4.63 ;
        RECT 18.25 4.13 18.35 4.23 ;
        RECT 18.25 3.73 18.35 3.83 ;
        RECT 18.45 27.33 18.55 27.43 ;
        RECT 18.45 26.93 18.55 27.03 ;
        RECT 18.45 26.53 18.55 26.63 ;
        RECT 18.45 26.13 18.55 26.23 ;
        RECT 18.45 25.73 18.55 25.83 ;
        RECT 18.45 25.33 18.55 25.43 ;
        RECT 18.45 24.93 18.55 25.03 ;
        RECT 18.45 24.53 18.55 24.63 ;
        RECT 18.45 24.13 18.55 24.23 ;
        RECT 18.45 23.73 18.55 23.83 ;
        RECT 18.45 23.33 18.55 23.43 ;
        RECT 18.45 22.93 18.55 23.03 ;
        RECT 18.45 22.53 18.55 22.63 ;
        RECT 18.45 22.13 18.55 22.23 ;
        RECT 18.45 21.73 18.55 21.83 ;
        RECT 18.45 21.33 18.55 21.43 ;
        RECT 18.45 20.93 18.55 21.03 ;
        RECT 18.45 20.53 18.55 20.63 ;
        RECT 18.45 20.13 18.55 20.23 ;
        RECT 18.45 19.73 18.55 19.83 ;
        RECT 18.45 19.33 18.55 19.43 ;
        RECT 18.45 18.93 18.55 19.03 ;
        RECT 18.45 18.53 18.55 18.63 ;
        RECT 18.45 18.13 18.55 18.23 ;
        RECT 18.45 17.73 18.55 17.83 ;
        RECT 18.45 17.33 18.55 17.43 ;
        RECT 18.45 16.93 18.55 17.03 ;
        RECT 18.45 16.53 18.55 16.63 ;
        RECT 18.45 16.13 18.55 16.23 ;
        RECT 18.45 15.73 18.55 15.83 ;
        RECT 18.45 15.33 18.55 15.43 ;
        RECT 18.45 14.93 18.55 15.03 ;
        RECT 18.45 14.53 18.55 14.63 ;
        RECT 18.45 14.13 18.55 14.23 ;
        RECT 18.45 13.73 18.55 13.83 ;
        RECT 18.45 13.33 18.55 13.43 ;
        RECT 18.45 12.93 18.55 13.03 ;
        RECT 18.45 12.53 18.55 12.63 ;
        RECT 18.45 12.13 18.55 12.23 ;
        RECT 18.45 11.73 18.55 11.83 ;
        RECT 18.45 11.33 18.55 11.43 ;
        RECT 18.45 10.93 18.55 11.03 ;
        RECT 18.45 10.53 18.55 10.63 ;
        RECT 18.45 10.13 18.55 10.23 ;
        RECT 18.45 9.73 18.55 9.83 ;
        RECT 18.45 9.33 18.55 9.43 ;
        RECT 18.45 8.93 18.55 9.03 ;
        RECT 18.45 8.53 18.55 8.63 ;
        RECT 18.45 8.13 18.55 8.23 ;
        RECT 18.45 7.73 18.55 7.83 ;
        RECT 18.45 7.33 18.55 7.43 ;
        RECT 18.45 6.93 18.55 7.03 ;
        RECT 18.45 6.53 18.55 6.63 ;
        RECT 18.45 6.13 18.55 6.23 ;
        RECT 18.45 5.73 18.55 5.83 ;
        RECT 18.45 5.33 18.55 5.43 ;
        RECT 18.45 4.93 18.55 5.03 ;
        RECT 18.45 4.53 18.55 4.63 ;
        RECT 18.45 4.13 18.55 4.23 ;
        RECT 18.45 3.73 18.55 3.83 ;
        RECT 23.745 52.26 23.845 52.36 ;
        RECT 23.745 52.03 23.845 52.13 ;
        RECT 23.745 51.8 23.845 51.9 ;
        RECT 23.745 51.57 23.845 51.67 ;
        RECT 23.745 51.34 23.845 51.44 ;
        RECT 23.745 51.11 23.845 51.21 ;
        RECT 23.745 50.88 23.845 50.98 ;
        RECT 23.745 50.65 23.845 50.75 ;
        RECT 23.745 50.42 23.845 50.52 ;
        RECT 23.745 50.19 23.845 50.29 ;
        RECT 23.745 49.96 23.845 50.06 ;
        RECT 23.745 49.73 23.845 49.83 ;
        RECT 23.95 27.33 24.05 27.43 ;
        RECT 23.95 26.93 24.05 27.03 ;
        RECT 23.95 26.53 24.05 26.63 ;
        RECT 23.95 26.13 24.05 26.23 ;
        RECT 23.95 25.73 24.05 25.83 ;
        RECT 23.95 25.33 24.05 25.43 ;
        RECT 23.95 24.93 24.05 25.03 ;
        RECT 23.95 24.53 24.05 24.63 ;
        RECT 23.95 24.13 24.05 24.23 ;
        RECT 23.95 23.73 24.05 23.83 ;
        RECT 23.95 23.33 24.05 23.43 ;
        RECT 23.95 22.93 24.05 23.03 ;
        RECT 23.95 22.53 24.05 22.63 ;
        RECT 23.95 22.13 24.05 22.23 ;
        RECT 23.95 21.73 24.05 21.83 ;
        RECT 23.95 21.33 24.05 21.43 ;
        RECT 23.95 20.93 24.05 21.03 ;
        RECT 23.95 20.53 24.05 20.63 ;
        RECT 23.95 20.13 24.05 20.23 ;
        RECT 23.95 19.73 24.05 19.83 ;
        RECT 23.95 19.33 24.05 19.43 ;
        RECT 23.95 18.93 24.05 19.03 ;
        RECT 23.95 18.53 24.05 18.63 ;
        RECT 23.95 18.13 24.05 18.23 ;
        RECT 23.95 17.73 24.05 17.83 ;
        RECT 23.95 17.33 24.05 17.43 ;
        RECT 23.95 16.93 24.05 17.03 ;
        RECT 23.95 16.53 24.05 16.63 ;
        RECT 23.95 16.13 24.05 16.23 ;
        RECT 23.95 15.73 24.05 15.83 ;
        RECT 23.95 15.33 24.05 15.43 ;
        RECT 23.95 14.93 24.05 15.03 ;
        RECT 23.95 14.53 24.05 14.63 ;
        RECT 23.95 14.13 24.05 14.23 ;
        RECT 23.95 13.73 24.05 13.83 ;
        RECT 23.95 13.33 24.05 13.43 ;
        RECT 23.95 12.93 24.05 13.03 ;
        RECT 23.95 12.53 24.05 12.63 ;
        RECT 23.95 12.13 24.05 12.23 ;
        RECT 23.95 11.73 24.05 11.83 ;
        RECT 23.95 11.33 24.05 11.43 ;
        RECT 23.95 10.93 24.05 11.03 ;
        RECT 23.95 10.53 24.05 10.63 ;
        RECT 23.95 10.13 24.05 10.23 ;
        RECT 23.95 9.73 24.05 9.83 ;
        RECT 23.95 9.33 24.05 9.43 ;
        RECT 23.95 8.93 24.05 9.03 ;
        RECT 23.95 8.53 24.05 8.63 ;
        RECT 23.95 8.13 24.05 8.23 ;
        RECT 23.95 7.73 24.05 7.83 ;
        RECT 23.95 7.33 24.05 7.43 ;
        RECT 23.95 6.93 24.05 7.03 ;
        RECT 23.95 6.53 24.05 6.63 ;
        RECT 23.95 6.13 24.05 6.23 ;
        RECT 23.95 5.73 24.05 5.83 ;
        RECT 23.95 5.33 24.05 5.43 ;
        RECT 23.95 4.93 24.05 5.03 ;
        RECT 23.95 4.53 24.05 4.63 ;
        RECT 23.95 4.13 24.05 4.23 ;
        RECT 23.95 3.73 24.05 3.83 ;
        RECT 23.975 52.26 24.075 52.36 ;
        RECT 23.975 52.03 24.075 52.13 ;
        RECT 23.975 51.8 24.075 51.9 ;
        RECT 23.975 51.57 24.075 51.67 ;
        RECT 23.975 51.34 24.075 51.44 ;
        RECT 23.975 51.11 24.075 51.21 ;
        RECT 23.975 50.88 24.075 50.98 ;
        RECT 23.975 50.65 24.075 50.75 ;
        RECT 23.975 50.42 24.075 50.52 ;
        RECT 23.975 50.19 24.075 50.29 ;
        RECT 23.975 49.96 24.075 50.06 ;
        RECT 23.975 49.73 24.075 49.83 ;
        RECT 24.15 27.33 24.25 27.43 ;
        RECT 24.15 26.93 24.25 27.03 ;
        RECT 24.15 26.53 24.25 26.63 ;
        RECT 24.15 26.13 24.25 26.23 ;
        RECT 24.15 25.73 24.25 25.83 ;
        RECT 24.15 25.33 24.25 25.43 ;
        RECT 24.15 24.93 24.25 25.03 ;
        RECT 24.15 24.53 24.25 24.63 ;
        RECT 24.15 24.13 24.25 24.23 ;
        RECT 24.15 23.73 24.25 23.83 ;
        RECT 24.15 23.33 24.25 23.43 ;
        RECT 24.15 22.93 24.25 23.03 ;
        RECT 24.15 22.53 24.25 22.63 ;
        RECT 24.15 22.13 24.25 22.23 ;
        RECT 24.15 21.73 24.25 21.83 ;
        RECT 24.15 21.33 24.25 21.43 ;
        RECT 24.15 20.93 24.25 21.03 ;
        RECT 24.15 20.53 24.25 20.63 ;
        RECT 24.15 20.13 24.25 20.23 ;
        RECT 24.15 19.73 24.25 19.83 ;
        RECT 24.15 19.33 24.25 19.43 ;
        RECT 24.15 18.93 24.25 19.03 ;
        RECT 24.15 18.53 24.25 18.63 ;
        RECT 24.15 18.13 24.25 18.23 ;
        RECT 24.15 17.73 24.25 17.83 ;
        RECT 24.15 17.33 24.25 17.43 ;
        RECT 24.15 16.93 24.25 17.03 ;
        RECT 24.15 16.53 24.25 16.63 ;
        RECT 24.15 16.13 24.25 16.23 ;
        RECT 24.15 15.73 24.25 15.83 ;
        RECT 24.15 15.33 24.25 15.43 ;
        RECT 24.15 14.93 24.25 15.03 ;
        RECT 24.15 14.53 24.25 14.63 ;
        RECT 24.15 14.13 24.25 14.23 ;
        RECT 24.15 13.73 24.25 13.83 ;
        RECT 24.15 13.33 24.25 13.43 ;
        RECT 24.15 12.93 24.25 13.03 ;
        RECT 24.15 12.53 24.25 12.63 ;
        RECT 24.15 12.13 24.25 12.23 ;
        RECT 24.15 11.73 24.25 11.83 ;
        RECT 24.15 11.33 24.25 11.43 ;
        RECT 24.15 10.93 24.25 11.03 ;
        RECT 24.15 10.53 24.25 10.63 ;
        RECT 24.15 10.13 24.25 10.23 ;
        RECT 24.15 9.73 24.25 9.83 ;
        RECT 24.15 9.33 24.25 9.43 ;
        RECT 24.15 8.93 24.25 9.03 ;
        RECT 24.15 8.53 24.25 8.63 ;
        RECT 24.15 8.13 24.25 8.23 ;
        RECT 24.15 7.73 24.25 7.83 ;
        RECT 24.15 7.33 24.25 7.43 ;
        RECT 24.15 6.93 24.25 7.03 ;
        RECT 24.15 6.53 24.25 6.63 ;
        RECT 24.15 6.13 24.25 6.23 ;
        RECT 24.15 5.73 24.25 5.83 ;
        RECT 24.15 5.33 24.25 5.43 ;
        RECT 24.15 4.93 24.25 5.03 ;
        RECT 24.15 4.53 24.25 4.63 ;
        RECT 24.15 4.13 24.25 4.23 ;
        RECT 24.15 3.73 24.25 3.83 ;
        RECT 24.205 52.26 24.305 52.36 ;
        RECT 24.205 52.03 24.305 52.13 ;
        RECT 24.205 51.8 24.305 51.9 ;
        RECT 24.205 51.57 24.305 51.67 ;
        RECT 24.205 51.34 24.305 51.44 ;
        RECT 24.205 51.11 24.305 51.21 ;
        RECT 24.205 50.88 24.305 50.98 ;
        RECT 24.205 50.65 24.305 50.75 ;
        RECT 24.205 50.42 24.305 50.52 ;
        RECT 24.205 50.19 24.305 50.29 ;
        RECT 24.205 49.96 24.305 50.06 ;
        RECT 24.205 49.73 24.305 49.83 ;
        RECT 24.35 27.33 24.45 27.43 ;
        RECT 24.35 26.93 24.45 27.03 ;
        RECT 24.35 26.53 24.45 26.63 ;
        RECT 24.35 26.13 24.45 26.23 ;
        RECT 24.35 25.73 24.45 25.83 ;
        RECT 24.35 25.33 24.45 25.43 ;
        RECT 24.35 24.93 24.45 25.03 ;
        RECT 24.35 24.53 24.45 24.63 ;
        RECT 24.35 24.13 24.45 24.23 ;
        RECT 24.35 23.73 24.45 23.83 ;
        RECT 24.35 23.33 24.45 23.43 ;
        RECT 24.35 22.93 24.45 23.03 ;
        RECT 24.35 22.53 24.45 22.63 ;
        RECT 24.35 22.13 24.45 22.23 ;
        RECT 24.35 21.73 24.45 21.83 ;
        RECT 24.35 21.33 24.45 21.43 ;
        RECT 24.35 20.93 24.45 21.03 ;
        RECT 24.35 20.53 24.45 20.63 ;
        RECT 24.35 20.13 24.45 20.23 ;
        RECT 24.35 19.73 24.45 19.83 ;
        RECT 24.35 19.33 24.45 19.43 ;
        RECT 24.35 18.93 24.45 19.03 ;
        RECT 24.35 18.53 24.45 18.63 ;
        RECT 24.35 18.13 24.45 18.23 ;
        RECT 24.35 17.73 24.45 17.83 ;
        RECT 24.35 17.33 24.45 17.43 ;
        RECT 24.35 16.93 24.45 17.03 ;
        RECT 24.35 16.53 24.45 16.63 ;
        RECT 24.35 16.13 24.45 16.23 ;
        RECT 24.35 15.73 24.45 15.83 ;
        RECT 24.35 15.33 24.45 15.43 ;
        RECT 24.35 14.93 24.45 15.03 ;
        RECT 24.35 14.53 24.45 14.63 ;
        RECT 24.35 14.13 24.45 14.23 ;
        RECT 24.35 13.73 24.45 13.83 ;
        RECT 24.35 13.33 24.45 13.43 ;
        RECT 24.35 12.93 24.45 13.03 ;
        RECT 24.35 12.53 24.45 12.63 ;
        RECT 24.35 12.13 24.45 12.23 ;
        RECT 24.35 11.73 24.45 11.83 ;
        RECT 24.35 11.33 24.45 11.43 ;
        RECT 24.35 10.93 24.45 11.03 ;
        RECT 24.35 10.53 24.45 10.63 ;
        RECT 24.35 10.13 24.45 10.23 ;
        RECT 24.35 9.73 24.45 9.83 ;
        RECT 24.35 9.33 24.45 9.43 ;
        RECT 24.35 8.93 24.45 9.03 ;
        RECT 24.35 8.53 24.45 8.63 ;
        RECT 24.35 8.13 24.45 8.23 ;
        RECT 24.35 7.73 24.45 7.83 ;
        RECT 24.35 7.33 24.45 7.43 ;
        RECT 24.35 6.93 24.45 7.03 ;
        RECT 24.35 6.53 24.45 6.63 ;
        RECT 24.35 6.13 24.45 6.23 ;
        RECT 24.35 5.73 24.45 5.83 ;
        RECT 24.35 5.33 24.45 5.43 ;
        RECT 24.35 4.93 24.45 5.03 ;
        RECT 24.35 4.53 24.45 4.63 ;
        RECT 24.35 4.13 24.45 4.23 ;
        RECT 24.35 3.73 24.45 3.83 ;
        RECT 24.435 52.26 24.535 52.36 ;
        RECT 24.435 52.03 24.535 52.13 ;
        RECT 24.435 51.8 24.535 51.9 ;
        RECT 24.435 51.57 24.535 51.67 ;
        RECT 24.435 51.34 24.535 51.44 ;
        RECT 24.435 51.11 24.535 51.21 ;
        RECT 24.435 50.88 24.535 50.98 ;
        RECT 24.435 50.65 24.535 50.75 ;
        RECT 24.435 50.42 24.535 50.52 ;
        RECT 24.435 50.19 24.535 50.29 ;
        RECT 24.435 49.96 24.535 50.06 ;
        RECT 24.435 49.73 24.535 49.83 ;
        RECT 24.665 52.26 24.765 52.36 ;
        RECT 24.665 52.03 24.765 52.13 ;
        RECT 24.665 51.8 24.765 51.9 ;
        RECT 24.665 51.57 24.765 51.67 ;
        RECT 24.665 51.34 24.765 51.44 ;
        RECT 24.665 51.11 24.765 51.21 ;
        RECT 24.665 50.88 24.765 50.98 ;
        RECT 24.665 50.65 24.765 50.75 ;
        RECT 24.665 50.42 24.765 50.52 ;
        RECT 24.665 50.19 24.765 50.29 ;
        RECT 24.665 49.96 24.765 50.06 ;
        RECT 24.665 49.73 24.765 49.83 ;
        RECT 24.895 52.26 24.995 52.36 ;
        RECT 24.895 52.03 24.995 52.13 ;
        RECT 24.895 51.8 24.995 51.9 ;
        RECT 24.895 51.57 24.995 51.67 ;
        RECT 24.895 51.34 24.995 51.44 ;
        RECT 24.895 51.11 24.995 51.21 ;
        RECT 24.895 50.88 24.995 50.98 ;
        RECT 24.895 50.65 24.995 50.75 ;
        RECT 24.895 50.42 24.995 50.52 ;
        RECT 24.895 50.19 24.995 50.29 ;
        RECT 24.895 49.96 24.995 50.06 ;
        RECT 24.895 49.73 24.995 49.83 ;
        RECT 25.125 52.26 25.225 52.36 ;
        RECT 25.125 52.03 25.225 52.13 ;
        RECT 25.125 51.8 25.225 51.9 ;
        RECT 25.125 51.57 25.225 51.67 ;
        RECT 25.125 51.34 25.225 51.44 ;
        RECT 25.125 51.11 25.225 51.21 ;
        RECT 25.125 50.88 25.225 50.98 ;
        RECT 25.125 50.65 25.225 50.75 ;
        RECT 25.125 50.42 25.225 50.52 ;
        RECT 25.125 50.19 25.225 50.29 ;
        RECT 25.125 49.96 25.225 50.06 ;
        RECT 25.125 49.73 25.225 49.83 ;
        RECT 25.355 52.26 25.455 52.36 ;
        RECT 25.355 52.03 25.455 52.13 ;
        RECT 25.355 51.8 25.455 51.9 ;
        RECT 25.355 51.57 25.455 51.67 ;
        RECT 25.355 51.34 25.455 51.44 ;
        RECT 25.355 51.11 25.455 51.21 ;
        RECT 25.355 50.88 25.455 50.98 ;
        RECT 25.355 50.65 25.455 50.75 ;
        RECT 25.355 50.42 25.455 50.52 ;
        RECT 25.355 50.19 25.455 50.29 ;
        RECT 25.355 49.96 25.455 50.06 ;
        RECT 25.355 49.73 25.455 49.83 ;
        RECT 25.585 52.26 25.685 52.36 ;
        RECT 25.585 52.03 25.685 52.13 ;
        RECT 25.585 51.8 25.685 51.9 ;
        RECT 25.585 51.57 25.685 51.67 ;
        RECT 25.585 51.34 25.685 51.44 ;
        RECT 25.585 51.11 25.685 51.21 ;
        RECT 25.585 50.88 25.685 50.98 ;
        RECT 25.585 50.65 25.685 50.75 ;
        RECT 25.585 50.42 25.685 50.52 ;
        RECT 25.585 50.19 25.685 50.29 ;
        RECT 25.585 49.96 25.685 50.06 ;
        RECT 25.585 49.73 25.685 49.83 ;
        RECT 25.815 52.26 25.915 52.36 ;
        RECT 25.815 52.03 25.915 52.13 ;
        RECT 25.815 51.8 25.915 51.9 ;
        RECT 25.815 51.57 25.915 51.67 ;
        RECT 25.815 51.34 25.915 51.44 ;
        RECT 25.815 51.11 25.915 51.21 ;
        RECT 25.815 50.88 25.915 50.98 ;
        RECT 25.815 50.65 25.915 50.75 ;
        RECT 25.815 50.42 25.915 50.52 ;
        RECT 25.815 50.19 25.915 50.29 ;
        RECT 25.815 49.96 25.915 50.06 ;
        RECT 25.815 49.73 25.915 49.83 ;
        RECT 26.045 52.26 26.145 52.36 ;
        RECT 26.045 52.03 26.145 52.13 ;
        RECT 26.045 51.8 26.145 51.9 ;
        RECT 26.045 51.57 26.145 51.67 ;
        RECT 26.045 51.34 26.145 51.44 ;
        RECT 26.045 51.11 26.145 51.21 ;
        RECT 26.045 50.88 26.145 50.98 ;
        RECT 26.045 50.65 26.145 50.75 ;
        RECT 26.045 50.42 26.145 50.52 ;
        RECT 26.045 50.19 26.145 50.29 ;
        RECT 26.045 49.96 26.145 50.06 ;
        RECT 26.045 49.73 26.145 49.83 ;
        RECT 26.275 52.26 26.375 52.36 ;
        RECT 26.275 52.03 26.375 52.13 ;
        RECT 26.275 51.8 26.375 51.9 ;
        RECT 26.275 51.57 26.375 51.67 ;
        RECT 26.275 51.34 26.375 51.44 ;
        RECT 26.275 51.11 26.375 51.21 ;
        RECT 26.275 50.88 26.375 50.98 ;
        RECT 26.275 50.65 26.375 50.75 ;
        RECT 26.275 50.42 26.375 50.52 ;
        RECT 26.275 50.19 26.375 50.29 ;
        RECT 26.275 49.96 26.375 50.06 ;
        RECT 26.275 49.73 26.375 49.83 ;
      LAYER M1 ;
        RECT 45 49.5 48 74.7 ;
        RECT 44.95 49.5 48 74.675 ;
        RECT 44.9 49.5 48 74.625 ;
        RECT 44.85 49.5 48 74.575 ;
        RECT 44.8 49.5 48 74.525 ;
        RECT 44.75 49.5 48 74.475 ;
        RECT 44.7 49.5 48 74.425 ;
        RECT 44.65 49.5 48 74.375 ;
        RECT 44.6 49.5 48 74.325 ;
        RECT 44.55 49.5 48 74.275 ;
        RECT 44.5 49.5 48 74.225 ;
        RECT 44.45 62 48 74.175 ;
        RECT 28.3 55 48 58 ;
        RECT 21.3 49.5 48 51 ;
        RECT 44.4 62 48 74.125 ;
        RECT 44.35 62 48 74.075 ;
        RECT 44.3 62 48 74.025 ;
        RECT 44.25 62 48 73.975 ;
        RECT 44.2 62 48 73.925 ;
        RECT 44.15 62 48 73.875 ;
        RECT 44.1 62 48 73.825 ;
        RECT 44.05 62 48 73.775 ;
        RECT 44 62 48 73.725 ;
        RECT 43.95 62 48 73.675 ;
        RECT 43.9 62 48 73.625 ;
        RECT 43.85 62 48 73.575 ;
        RECT 43.8 62 48 73.525 ;
        RECT 43.75 62 48 73.475 ;
        RECT 43.7 62 48 73.425 ;
        RECT 43.65 62 48 73.375 ;
        RECT 43.6 62 48 73.325 ;
        RECT 43.55 62 48 73.275 ;
        RECT 43.5 62 48 73.225 ;
        RECT 43.45 62 48 73.175 ;
        RECT 43.4 62 48 73.125 ;
        RECT 43.35 62 48 73.075 ;
        RECT 43.3 62 48 73.025 ;
        RECT 43.25 62 48 72.975 ;
        RECT 43.2 62 48 72.925 ;
        RECT 43.15 62 48 72.875 ;
        RECT 43.1 62 48 72.825 ;
        RECT 43.05 62 48 72.775 ;
        RECT 43 62 48 72.725 ;
        RECT 42.95 62 48 72.675 ;
        RECT 42.9 62 48 72.625 ;
        RECT 42.85 62 48 72.575 ;
        RECT 42.8 62 48 72.525 ;
        RECT 42.75 62 48 72.475 ;
        RECT 42.7 62 48 72.425 ;
        RECT 42.65 62 48 72.375 ;
        RECT 42.6 62 48 72.325 ;
        RECT 42.55 62 48 72.275 ;
        RECT 42.5 62 48 72.225 ;
        RECT 42.45 62 48 72.175 ;
        RECT 42.4 62 48 72.125 ;
        RECT 42.35 62 48 72.075 ;
        RECT 42.3 62 48 72.025 ;
        RECT 42.25 62 48 71.975 ;
        RECT 42.2 62 48 71.925 ;
        RECT 42.15 62 48 71.875 ;
        RECT 42.1 62 48 71.825 ;
        RECT 42.05 62 48 71.775 ;
        RECT 42 62 48 71.725 ;
        RECT 41.95 62 48 71.675 ;
        RECT 41.9 62 48 71.625 ;
        RECT 41.85 62 48 71.575 ;
        RECT 41.8 62 48 71.525 ;
        RECT 41.75 62 48 71.475 ;
        RECT 41.7 62 48 71.425 ;
        RECT 41.65 62 48 71.375 ;
        RECT 41.6 62 48 71.325 ;
        RECT 41.55 62 48 71.275 ;
        RECT 41.5 62 48 71.225 ;
        RECT 41.45 62 48 71.175 ;
        RECT 41.4 62 48 71.125 ;
        RECT 41.35 62 48 71.075 ;
        RECT 41.3 62 48 71.025 ;
        RECT 41.25 62 48 70.975 ;
        RECT 41.2 62 48 70.925 ;
        RECT 41.15 62 48 70.875 ;
        RECT 41.1 62 48 70.825 ;
        RECT 41.05 62 48 70.775 ;
        RECT 41 62 48 70.725 ;
        RECT 40.95 62 48 70.675 ;
        RECT 40.9 62 48 70.625 ;
        RECT 40.85 62 48 70.575 ;
        RECT 40.8 62 48 70.525 ;
        RECT 40.75 62 48 70.475 ;
        RECT 40.7 62 48 70.425 ;
        RECT 40.65 62 48 70.375 ;
        RECT 40.6 62 48 70.325 ;
        RECT 40.55 62 48 70.275 ;
        RECT 40.5 62 48 70.225 ;
        RECT 32.3 55 40.5 62.025 ;
        RECT 37.5 49.5 40.5 67.225 ;
        RECT 40.45 62 48 70.175 ;
        RECT 40.4 62 48 70.125 ;
        RECT 40.35 62 48 70.075 ;
        RECT 40.3 62 48 70.025 ;
        RECT 40.25 62 48 69.975 ;
        RECT 40.2 62 48 69.925 ;
        RECT 40.15 62 48 69.875 ;
        RECT 40.1 62 48 69.825 ;
        RECT 40.05 62 48 69.775 ;
        RECT 40 62 48 69.725 ;
        RECT 39.95 62 48 69.675 ;
        RECT 39.9 62 48 69.625 ;
        RECT 39.85 62 48 69.575 ;
        RECT 39.8 62 48 69.525 ;
        RECT 39.75 62 48 69.475 ;
        RECT 39.7 62 48 69.425 ;
        RECT 39.65 62 48 69.375 ;
        RECT 39.6 62 48 69.325 ;
        RECT 39.55 62 48 69.275 ;
        RECT 39.5 62 48 69.225 ;
        RECT 39.45 62 48 69.175 ;
        RECT 39.4 62 48 69.125 ;
        RECT 39.35 62 48 69.075 ;
        RECT 39.3 62 48 69.025 ;
        RECT 39.25 62 48 68.975 ;
        RECT 39.2 62 48 68.925 ;
        RECT 39.15 62 48 68.875 ;
        RECT 39.1 62 48 68.825 ;
        RECT 39.05 62 48 68.775 ;
        RECT 39 62 48 68.725 ;
        RECT 38.95 62 48 68.675 ;
        RECT 38.9 62 48 68.625 ;
        RECT 38.85 62 48 68.575 ;
        RECT 38.8 62 48 68.525 ;
        RECT 38.75 62 48 68.475 ;
        RECT 38.7 62 48 68.425 ;
        RECT 38.65 62 48 68.375 ;
        RECT 38.6 62 48 68.325 ;
        RECT 38.55 62 48 68.275 ;
        RECT 38.5 62 48 68.225 ;
        RECT 38.45 62 48 68.175 ;
        RECT 38.4 62 48 68.125 ;
        RECT 38.35 62 48 68.075 ;
        RECT 38.3 62 48 68.025 ;
        RECT 38.25 62 48 67.975 ;
        RECT 38.2 62 48 67.925 ;
        RECT 38.15 62 48 67.875 ;
        RECT 38.1 62 48 67.825 ;
        RECT 38.05 62 48 67.775 ;
        RECT 38 62 48 67.725 ;
        RECT 37.95 62 48 67.675 ;
        RECT 37.9 62 48 67.625 ;
        RECT 37.85 62 48 67.575 ;
        RECT 37.8 62 48 67.525 ;
        RECT 37.75 62 48 67.475 ;
        RECT 37.7 62 48 67.425 ;
        RECT 37.65 62 48 67.375 ;
        RECT 37.6 62 48 67.325 ;
        RECT 37.55 62 48 67.275 ;
        RECT 37.45 62 48 67.175 ;
        RECT 37.4 62 48 67.125 ;
        RECT 37.35 62 48 67.075 ;
        RECT 37.3 62 48 67.025 ;
        RECT 37.25 62 48 66.975 ;
        RECT 37.2 62 48 66.925 ;
        RECT 37.15 62 48 66.875 ;
        RECT 37.1 62 48 66.825 ;
        RECT 37.05 62 48 66.775 ;
        RECT 37 62 48 66.725 ;
        RECT 19.8 49.475 37 49.525 ;
        RECT 36.95 62 48 66.675 ;
        RECT 19.75 49.425 36.95 49.475 ;
        RECT 36.9 62 48 66.625 ;
        RECT 19.7 49.375 36.9 49.425 ;
        RECT 36.85 62 48 66.575 ;
        RECT 19.65 49.325 36.85 49.375 ;
        RECT 36.8 62 48 66.525 ;
        RECT 19.6 49.275 36.8 49.325 ;
        RECT 36.75 62 48 66.475 ;
        RECT 19.55 49.225 36.75 49.275 ;
        RECT 36.7 62 48 66.425 ;
        RECT 19.5 49.175 36.7 49.225 ;
        RECT 36.65 62 48 66.375 ;
        RECT 19.45 49.125 36.65 49.175 ;
        RECT 36.6 62 48 66.325 ;
        RECT 19.4 49.075 36.6 49.125 ;
        RECT 36.55 62 48 66.275 ;
        RECT 19.35 49.025 36.55 49.075 ;
        RECT 36.5 62 48 66.225 ;
        RECT 19.3 48.975 36.5 49.025 ;
        RECT 36.45 62 48 66.175 ;
        RECT 19.25 48.925 36.45 48.975 ;
        RECT 36.4 62 48 66.125 ;
        RECT 19.2 48.875 36.4 48.925 ;
        RECT 36.35 62 48 66.075 ;
        RECT 19.15 48.825 36.35 48.875 ;
        RECT 36.3 62 48 66.025 ;
        RECT 19.1 48.775 36.3 48.825 ;
        RECT 36.25 62 48 65.975 ;
        RECT 19.05 48.725 36.25 48.775 ;
        RECT 36.2 62 48 65.925 ;
        RECT 19 48.675 36.2 48.725 ;
        RECT 36.15 62 48 65.875 ;
        RECT 18.95 48.625 36.15 48.675 ;
        RECT 36.1 62 48 65.825 ;
        RECT 18.9 48.575 36.1 48.625 ;
        RECT 36.05 62 48 65.775 ;
        RECT 18.85 48.525 36.05 48.575 ;
        RECT 36 62 48 65.725 ;
        RECT 18.8 48.475 36 48.525 ;
        RECT 35.95 62 48 65.675 ;
        RECT 18.75 48.425 35.95 48.475 ;
        RECT 35.9 62 48 65.625 ;
        RECT 18.7 48.375 35.9 48.425 ;
        RECT 35.85 62 48 65.575 ;
        RECT 18.65 48.325 35.85 48.375 ;
        RECT 35.8 62 48 65.525 ;
        RECT 18.6 48.275 35.8 48.325 ;
        RECT 35.75 62 48 65.475 ;
        RECT 18.55 48.225 35.75 48.275 ;
        RECT 35.7 62 48 65.425 ;
        RECT 18.5 48.175 35.7 48.225 ;
        RECT 35.65 62 48 65.375 ;
        RECT 18.45 48.125 35.65 48.175 ;
        RECT 35.6 62 48 65.325 ;
        RECT 18.4 48.075 35.6 48.125 ;
        RECT 35.55 62 48 65.275 ;
        RECT 18.35 48.025 35.55 48.075 ;
        RECT 35.5 62 48 65.225 ;
        RECT 32 47.975 35.5 51 ;
        RECT 35.45 62 48 65.175 ;
        RECT 32 47.925 35.45 51 ;
        RECT 35.4 62 48 65.125 ;
        RECT 32 47.875 35.4 51 ;
        RECT 35.35 62 48 65.075 ;
        RECT 32 47.825 35.35 51 ;
        RECT 35.3 62 48 65.025 ;
        RECT 32 47.775 35.3 51 ;
        RECT 35.25 62 48 64.975 ;
        RECT 32 47.725 35.25 51 ;
        RECT 35.2 62 48 64.925 ;
        RECT 32 47.675 35.2 51 ;
        RECT 35.15 62 48 64.875 ;
        RECT 32 47.625 35.15 51 ;
        RECT 35.1 62 48 64.825 ;
        RECT 32 47.575 35.1 51 ;
        RECT 35.05 62 48 64.775 ;
        RECT 32 47.525 35.05 51 ;
        RECT 35 62 48 64.725 ;
        RECT 32 47.475 35 51 ;
        RECT 34.95 62 48 64.675 ;
        RECT 32 47.425 34.95 51 ;
        RECT 34.9 62 48 64.625 ;
        RECT 32 47.375 34.9 51 ;
        RECT 34.85 62 48 64.575 ;
        RECT 32 47.325 34.85 51 ;
        RECT 34.8 62 48 64.525 ;
        RECT 32 47.275 34.8 51 ;
        RECT 34.75 62 48 64.475 ;
        RECT 32 47.225 34.75 51 ;
        RECT 34.7 62 48 64.425 ;
        RECT 32 47.175 34.7 51 ;
        RECT 34.65 62 48 64.375 ;
        RECT 32 47.125 34.65 51 ;
        RECT 34.6 62 48 64.325 ;
        RECT 32 47.075 34.6 51 ;
        RECT 34.55 62 48 64.275 ;
        RECT 32 47.025 34.55 51 ;
        RECT 34.5 62 48 64.225 ;
        RECT 32 46.975 34.5 51 ;
        RECT 34.45 62 48 64.175 ;
        RECT 32 46.925 34.45 51 ;
        RECT 34.4 62 48 64.125 ;
        RECT 32 46.875 34.4 51 ;
        RECT 34.35 62 48 64.075 ;
        RECT 32 46.825 34.35 51 ;
        RECT 34.3 62 48 64.025 ;
        RECT 32 46.775 34.3 51 ;
        RECT 34.25 62 48 63.975 ;
        RECT 32 46.725 34.25 51 ;
        RECT 34.2 62 48 63.925 ;
        RECT 32 46.675 34.2 51 ;
        RECT 34.15 62 48 63.875 ;
        RECT 32 46.625 34.15 51 ;
        RECT 34.1 62 48 63.825 ;
        RECT 32 46.575 34.1 51 ;
        RECT 34.05 62 48 63.775 ;
        RECT 32 46.525 34.05 51 ;
        RECT 34 62 48 63.725 ;
        RECT 32 46.475 34 51 ;
        RECT 33.95 62 48 63.675 ;
        RECT 32 46.425 33.95 51 ;
        RECT 33.9 62 48 63.625 ;
        RECT 32 46.375 33.9 51 ;
        RECT 33.85 62 48 63.575 ;
        RECT 32 46.325 33.85 51 ;
        RECT 33.8 62 48 63.525 ;
        RECT 32 46.275 33.8 51 ;
        RECT 33.75 62 48 63.475 ;
        RECT 32 46.225 33.75 51 ;
        RECT 33.7 62 48 63.425 ;
        RECT 32 46.175 33.7 51 ;
        RECT 33.65 62 48 63.375 ;
        RECT 32 46.125 33.65 51 ;
        RECT 33.6 62 48 63.325 ;
        RECT 32 46.075 33.6 51 ;
        RECT 33.55 62 48 63.275 ;
        RECT 32 46.025 33.55 51 ;
        RECT 33.5 62 48 63.225 ;
        RECT 25.3 48 33.5 55.025 ;
        RECT 32 42.5 33.5 61.725 ;
        RECT 33.45 62 48 63.175 ;
        RECT 33.4 62 48 63.125 ;
        RECT 33.35 62 48 63.075 ;
        RECT 33.3 62 48 63.025 ;
        RECT 33.25 62 48 62.975 ;
        RECT 33.2 62 48 62.925 ;
        RECT 33.15 62 48 62.875 ;
        RECT 33.1 62 48 62.825 ;
        RECT 33.05 62 48 62.775 ;
        RECT 33 62 48 62.725 ;
        RECT 32.95 62 48 62.675 ;
        RECT 32.9 62 48 62.625 ;
        RECT 32.85 62 48 62.575 ;
        RECT 32.8 62 48 62.525 ;
        RECT 32.75 62 48 62.475 ;
        RECT 32.7 62 48 62.425 ;
        RECT 32.65 62 48 62.375 ;
        RECT 32.6 62 48 62.325 ;
        RECT 32.55 62 48 62.275 ;
        RECT 32.5 62 48 62.225 ;
        RECT 32.45 62 48 62.175 ;
        RECT 32.4 62 48 62.125 ;
        RECT 32.35 62 48 62.075 ;
        RECT 32.25 55 40.5 61.975 ;
        RECT 32.2 55 40.5 61.925 ;
        RECT 32.15 55 40.5 61.875 ;
        RECT 32.1 55 40.5 61.825 ;
        RECT 32.05 55 40.5 61.775 ;
        RECT 31.95 55 40.5 61.675 ;
        RECT 14.3 42.5 33.5 44 ;
        RECT 31.9 55 40.5 61.625 ;
        RECT 31.85 55 40.5 61.575 ;
        RECT 31.8 55 40.5 61.525 ;
        RECT 31.75 55 40.5 61.475 ;
        RECT 31.7 55 40.5 61.425 ;
        RECT 31.65 55 40.5 61.375 ;
        RECT 31.6 55 40.5 61.325 ;
        RECT 31.55 55 40.5 61.275 ;
        RECT 31.5 55 40.5 61.225 ;
        RECT 31.45 55 40.5 61.175 ;
        RECT 31.4 55 40.5 61.125 ;
        RECT 31.35 55 40.5 61.075 ;
        RECT 31.3 55 40.5 61.025 ;
        RECT 31.25 55 40.5 60.975 ;
        RECT 31.2 55 40.5 60.925 ;
        RECT 31.15 55 40.5 60.875 ;
        RECT 31.1 55 40.5 60.825 ;
        RECT 31.05 55 40.5 60.775 ;
        RECT 31 55 40.5 60.725 ;
        RECT 30.95 55 40.5 60.675 ;
        RECT 30.9 55 40.5 60.625 ;
        RECT 30.85 55 40.5 60.575 ;
        RECT 30.8 55 40.5 60.525 ;
        RECT 30.75 55 40.5 60.475 ;
        RECT 30.7 55 40.5 60.425 ;
        RECT 30.65 55 40.5 60.375 ;
        RECT 30.6 55 40.5 60.325 ;
        RECT 30.55 55 40.5 60.275 ;
        RECT 30.5 55 40.5 60.225 ;
        RECT 30.45 55 40.5 60.175 ;
        RECT 30.4 55 40.5 60.125 ;
        RECT 30.35 55 40.5 60.075 ;
        RECT 30.3 55 40.5 60.025 ;
        RECT 30.25 55 40.5 59.975 ;
        RECT 30.2 55 40.5 59.925 ;
        RECT 30.15 55 40.5 59.875 ;
        RECT 30.1 55 40.5 59.825 ;
        RECT 30.05 55 40.5 59.775 ;
        RECT 30 55 40.5 59.725 ;
        RECT 12.8 42.475 30 42.525 ;
        RECT 29.95 55 40.5 59.675 ;
        RECT 12.75 42.425 29.95 42.475 ;
        RECT 29.9 55 40.5 59.625 ;
        RECT 12.7 42.375 29.9 42.425 ;
        RECT 29.85 55 40.5 59.575 ;
        RECT 12.65 42.325 29.85 42.375 ;
        RECT 29.8 55 40.5 59.525 ;
        RECT 12.6 42.275 29.8 42.325 ;
        RECT 29.75 55 40.5 59.475 ;
        RECT 12.55 42.225 29.75 42.275 ;
        RECT 29.7 55 40.5 59.425 ;
        RECT 12.5 42.175 29.7 42.225 ;
        RECT 29.65 55 40.5 59.375 ;
        RECT 12.45 42.125 29.65 42.175 ;
        RECT 29.6 55 40.5 59.325 ;
        RECT 12.4 42.075 29.6 42.125 ;
        RECT 29.55 55 40.5 59.275 ;
        RECT 12.35 42.025 29.55 42.075 ;
        RECT 29.5 55 40.5 59.225 ;
        RECT 12.3 41.975 29.5 42.025 ;
        RECT 29.45 55 40.5 59.175 ;
        RECT 12.25 41.925 29.45 41.975 ;
        RECT 29.4 55 40.5 59.125 ;
        RECT 12.2 41.875 29.4 41.925 ;
        RECT 29.35 55 40.5 59.075 ;
        RECT 12.15 41.825 29.35 41.875 ;
        RECT 29.3 55 40.5 59.025 ;
        RECT 12.1 41.775 29.3 41.825 ;
        RECT 29.25 55 40.5 58.975 ;
        RECT 12.05 41.725 29.25 41.775 ;
        RECT 29.2 55 40.5 58.925 ;
        RECT 12 41.675 29.2 41.725 ;
        RECT 29.15 55 40.5 58.875 ;
        RECT 11.95 41.625 29.15 41.675 ;
        RECT 29.1 55 40.5 58.825 ;
        RECT 11.9 41.575 29.1 41.625 ;
        RECT 29.05 55 40.5 58.775 ;
        RECT 11.85 41.525 29.05 41.575 ;
        RECT 29 55 40.5 58.725 ;
        RECT 11.8 41.475 29 41.525 ;
        RECT 28.95 55 40.5 58.675 ;
        RECT 11.75 41.425 28.95 41.475 ;
        RECT 28.9 55 40.5 58.625 ;
        RECT 11.7 41.375 28.9 41.425 ;
        RECT 28.85 55 40.5 58.575 ;
        RECT 11.65 41.325 28.85 41.375 ;
        RECT 28.8 55 40.5 58.525 ;
        RECT 11.6 41.275 28.8 41.325 ;
        RECT 28.75 55 40.5 58.475 ;
        RECT 11.55 41.225 28.75 41.275 ;
        RECT 28.7 55 40.5 58.425 ;
        RECT 11.5 41.175 28.7 41.225 ;
        RECT 28.65 55 40.5 58.375 ;
        RECT 11.45 41.125 28.65 41.175 ;
        RECT 28.6 55 40.5 58.325 ;
        RECT 11.4 41.075 28.6 41.125 ;
        RECT 28.55 55 40.5 58.275 ;
        RECT 11.35 41.025 28.55 41.075 ;
        RECT 28.5 55 40.5 58.225 ;
        RECT 23.5 40.975 28.5 44 ;
        RECT 28.45 55 40.5 58.175 ;
        RECT 23.5 40.925 28.45 44 ;
        RECT 28.4 55 40.5 58.125 ;
        RECT 23.5 40.875 28.4 44 ;
        RECT 28.35 55 40.5 58.075 ;
        RECT 23.5 40.825 28.35 44 ;
        RECT 28.3 55 40.5 58.025 ;
        RECT 23.5 40.775 28.3 44 ;
        RECT 28.25 55 48 57.975 ;
        RECT 23.5 40.725 28.25 44 ;
        RECT 28.2 55 48 57.925 ;
        RECT 23.5 40.675 28.2 44 ;
        RECT 28.15 55 48 57.875 ;
        RECT 23.5 40.625 28.15 44 ;
        RECT 28.1 55 48 57.825 ;
        RECT 23.5 40.575 28.1 44 ;
        RECT 28.05 55 48 57.775 ;
        RECT 23.5 40.525 28.05 44 ;
        RECT 28 55 48 57.725 ;
        RECT 18.3 41 28 48.025 ;
        RECT 23.5 40.475 28 53.225 ;
        RECT 27.95 55 48 57.675 ;
        RECT 23.5 40.425 27.95 53.225 ;
        RECT 27.9 55 48 57.625 ;
        RECT 23.5 40.375 27.9 53.225 ;
        RECT 27.85 55 48 57.575 ;
        RECT 23.5 40.325 27.85 53.225 ;
        RECT 27.8 55 48 57.525 ;
        RECT 23.5 40.275 27.8 53.225 ;
        RECT 27.75 55 48 57.475 ;
        RECT 23.5 40.225 27.75 53.225 ;
        RECT 27.7 55 48 57.425 ;
        RECT 23.5 40.175 27.7 53.225 ;
        RECT 27.65 55 48 57.375 ;
        RECT 23.5 40.125 27.65 53.225 ;
        RECT 27.6 55 48 57.325 ;
        RECT 23.5 40.075 27.6 53.225 ;
        RECT 27.55 55 48 57.275 ;
        RECT 23.5 40.025 27.55 53.225 ;
        RECT 27.5 55 48 57.225 ;
        RECT 23.5 39.975 27.5 53.225 ;
        RECT 27.45 55 48 57.175 ;
        RECT 23.5 39.925 27.45 53.225 ;
        RECT 27.4 55 48 57.125 ;
        RECT 23.5 39.875 27.4 53.225 ;
        RECT 27.35 55 48 57.075 ;
        RECT 23.5 39.825 27.35 53.225 ;
        RECT 27.3 55 48 57.025 ;
        RECT 23.5 39.775 27.3 53.225 ;
        RECT 27.25 55 48 56.975 ;
        RECT 23.5 39.725 27.25 53.225 ;
        RECT 27.2 55 48 56.925 ;
        RECT 23.5 39.675 27.2 53.225 ;
        RECT 27.15 55 48 56.875 ;
        RECT 23.5 39.625 27.15 53.225 ;
        RECT 27.1 55 48 56.825 ;
        RECT 23.5 39.575 27.1 53.225 ;
        RECT 27.05 55 48 56.775 ;
        RECT 23.5 39.525 27.05 53.225 ;
        RECT 27 55 48 56.725 ;
        RECT 23.5 39.475 27 53.225 ;
        RECT 26.95 55 48 56.675 ;
        RECT 23.5 39.425 26.95 53.225 ;
        RECT 26.9 55 48 56.625 ;
        RECT 23.5 39.375 26.9 53.225 ;
        RECT 26.85 55 48 56.575 ;
        RECT 23.5 39.325 26.85 53.225 ;
        RECT 26.8 55 48 56.525 ;
        RECT 23.5 39.275 26.8 53.225 ;
        RECT 26.75 55 48 56.475 ;
        RECT 23.5 39.225 26.75 53.225 ;
        RECT 26.7 55 48 56.425 ;
        RECT 23.5 39.175 26.7 53.225 ;
        RECT 26.65 55 48 56.375 ;
        RECT 23.5 39.125 26.65 53.225 ;
        RECT 26.6 55 48 56.325 ;
        RECT 23.5 39.075 26.6 53.225 ;
        RECT 26.55 55 48 56.275 ;
        RECT 23.5 39.025 26.55 53.225 ;
        RECT 26.5 55 48 56.225 ;
        RECT 23.5 0 26.5 53.225 ;
        RECT 26.45 55 48 56.175 ;
        RECT 26.4 55 48 56.125 ;
        RECT 26.35 55 48 56.075 ;
        RECT 26.3 55 48 56.025 ;
        RECT 26.25 55 48 55.975 ;
        RECT 26.2 55 48 55.925 ;
        RECT 26.15 55 48 55.875 ;
        RECT 26.1 55 48 55.825 ;
        RECT 26.05 55 48 55.775 ;
        RECT 26 55 48 55.725 ;
        RECT 25.95 55 48 55.675 ;
        RECT 25.9 55 48 55.625 ;
        RECT 25.85 55 48 55.575 ;
        RECT 25.8 55 48 55.525 ;
        RECT 25.75 55 48 55.475 ;
        RECT 25.7 55 48 55.425 ;
        RECT 25.65 55 48 55.375 ;
        RECT 25.6 55 48 55.325 ;
        RECT 25.55 55 48 55.275 ;
        RECT 25.5 55 48 55.225 ;
        RECT 25.45 55 48 55.175 ;
        RECT 25.4 55 48 55.125 ;
        RECT 25.35 55 48 55.075 ;
        RECT 25.25 48 33.5 54.975 ;
        RECT 25.2 48 33.5 54.925 ;
        RECT 25.15 48 33.5 54.875 ;
        RECT 25.1 48 33.5 54.825 ;
        RECT 25.05 48 33.5 54.775 ;
        RECT 25 48 33.5 54.725 ;
        RECT 24.95 48 33.5 54.675 ;
        RECT 24.9 48 33.5 54.625 ;
        RECT 24.85 48 33.5 54.575 ;
        RECT 24.8 48 33.5 54.525 ;
        RECT 24.75 48 33.5 54.475 ;
        RECT 24.7 48 33.5 54.425 ;
        RECT 24.65 48 33.5 54.375 ;
        RECT 24.6 48 33.5 54.325 ;
        RECT 24.55 48 33.5 54.275 ;
        RECT 24.5 48 33.5 54.225 ;
        RECT 24.45 48 33.5 54.175 ;
        RECT 24.4 48 33.5 54.125 ;
        RECT 24.35 48 33.5 54.075 ;
        RECT 24.3 48 33.5 54.025 ;
        RECT 24.25 48 33.5 53.975 ;
        RECT 24.2 48 33.5 53.925 ;
        RECT 24.15 48 33.5 53.875 ;
        RECT 24.1 48 33.5 53.825 ;
        RECT 24.05 48 33.5 53.775 ;
        RECT 24 48 33.5 53.725 ;
        RECT 23.95 48 33.5 53.675 ;
        RECT 23.9 48 33.5 53.625 ;
        RECT 23.85 48 33.5 53.575 ;
        RECT 23.8 48 33.5 53.525 ;
        RECT 23.75 48 33.5 53.475 ;
        RECT 23.7 48 33.5 53.425 ;
        RECT 23.65 48 33.5 53.375 ;
        RECT 23.6 48 33.5 53.325 ;
        RECT 23.55 48 33.5 53.275 ;
        RECT 23.45 48 33.5 53.175 ;
        RECT 7.3 34 26.5 37 ;
        RECT 1.3 27 26.5 30 ;
        RECT 1.3 20 26.5 23 ;
        RECT 1.3 13 26.5 16 ;
        RECT 1.3 6 26.5 9 ;
        RECT 1.3 0 26.5 2 ;
        RECT 23.4 48 33.5 53.125 ;
        RECT 23.35 48 33.5 53.075 ;
        RECT 23.3 48 33.5 53.025 ;
        RECT 23.25 48 33.5 52.975 ;
        RECT 23.2 48 33.5 52.925 ;
        RECT 23.15 48 33.5 52.875 ;
        RECT 23.1 48 33.5 52.825 ;
        RECT 23.05 48 33.5 52.775 ;
        RECT 23 48 33.5 52.725 ;
        RECT 22.95 48 33.5 52.675 ;
        RECT 22.9 48 33.5 52.625 ;
        RECT 22.85 48 33.5 52.575 ;
        RECT 22.8 48 33.5 52.525 ;
        RECT 22.75 48 33.5 52.475 ;
        RECT 22.7 48 33.5 52.425 ;
        RECT 22.65 48 33.5 52.375 ;
        RECT 22.6 48 33.5 52.325 ;
        RECT 22.55 48 33.5 52.275 ;
        RECT 22.5 48 33.5 52.225 ;
        RECT 22.45 48 33.5 52.175 ;
        RECT 22.4 48 33.5 52.125 ;
        RECT 22.35 48 33.5 52.075 ;
        RECT 22.3 48 33.5 52.025 ;
        RECT 22.25 48 33.5 51.975 ;
        RECT 22.2 48 33.5 51.925 ;
        RECT 22.15 48 33.5 51.875 ;
        RECT 22.1 48 33.5 51.825 ;
        RECT 22.05 48 33.5 51.775 ;
        RECT 22 48 33.5 51.725 ;
        RECT 21.95 48 33.5 51.675 ;
        RECT 21.9 48 33.5 51.625 ;
        RECT 21.85 48 33.5 51.575 ;
        RECT 21.8 48 33.5 51.525 ;
        RECT 21.75 48 33.5 51.475 ;
        RECT 21.7 48 33.5 51.425 ;
        RECT 21.65 48 33.5 51.375 ;
        RECT 21.6 48 33.5 51.325 ;
        RECT 21.55 48 33.5 51.275 ;
        RECT 21.5 48 33.5 51.225 ;
        RECT 21.45 48 33.5 51.175 ;
        RECT 21.4 48 33.5 51.125 ;
        RECT 21.35 48 33.5 51.075 ;
        RECT 21.3 48 33.5 51.025 ;
        RECT 21.25 49.5 48 50.975 ;
        RECT 21.2 49.5 48 50.925 ;
        RECT 21.15 49.5 48 50.875 ;
        RECT 21.1 49.5 48 50.825 ;
        RECT 21.05 49.5 48 50.775 ;
        RECT 21 49.5 48 50.725 ;
        RECT 20.95 49.5 48 50.675 ;
        RECT 20.9 49.5 48 50.625 ;
        RECT 20.85 49.5 48 50.575 ;
        RECT 20.8 49.5 48 50.525 ;
        RECT 20.75 49.5 48 50.475 ;
        RECT 20.7 49.5 48 50.425 ;
        RECT 20.65 49.5 48 50.375 ;
        RECT 20.6 49.5 48 50.325 ;
        RECT 20.55 49.5 48 50.275 ;
        RECT 20.5 49.5 48 50.225 ;
        RECT 20.45 49.5 48 50.175 ;
        RECT 20.4 49.5 48 50.125 ;
        RECT 20.35 49.5 48 50.075 ;
        RECT 20.3 49.5 48 50.025 ;
        RECT 20.25 49.5 48 49.975 ;
        RECT 20.2 49.5 48 49.925 ;
        RECT 20.15 49.5 48 49.875 ;
        RECT 20.1 49.5 48 49.825 ;
        RECT 20.05 49.5 48 49.775 ;
        RECT 20 49.5 48 49.725 ;
        RECT 19.95 49.5 48 49.675 ;
        RECT 19.9 49.5 48 49.625 ;
        RECT 19.85 49.5 48 49.575 ;
        RECT 11.3 34 19.5 41.025 ;
        RECT 16.5 0 19.5 46.225 ;
        RECT 18.25 41 28 47.975 ;
        RECT 18.2 41 28 47.925 ;
        RECT 18.15 41 28 47.875 ;
        RECT 18.1 41 28 47.825 ;
        RECT 18.05 41 28 47.775 ;
        RECT 18 41 28 47.725 ;
        RECT 17.95 41 28 47.675 ;
        RECT 17.9 41 28 47.625 ;
        RECT 17.85 41 28 47.575 ;
        RECT 17.8 41 28 47.525 ;
        RECT 17.75 41 28 47.475 ;
        RECT 17.7 41 28 47.425 ;
        RECT 17.65 41 28 47.375 ;
        RECT 17.6 41 28 47.325 ;
        RECT 17.55 41 28 47.275 ;
        RECT 17.5 41 28 47.225 ;
        RECT 17.45 41 28 47.175 ;
        RECT 17.4 41 28 47.125 ;
        RECT 17.35 41 28 47.075 ;
        RECT 17.3 41 28 47.025 ;
        RECT 17.25 41 28 46.975 ;
        RECT 17.2 41 28 46.925 ;
        RECT 17.15 41 28 46.875 ;
        RECT 17.1 41 28 46.825 ;
        RECT 17.05 41 28 46.775 ;
        RECT 17 41 28 46.725 ;
        RECT 16.95 41 28 46.675 ;
        RECT 16.9 41 28 46.625 ;
        RECT 16.85 41 28 46.575 ;
        RECT 16.8 41 28 46.525 ;
        RECT 16.75 41 28 46.475 ;
        RECT 16.7 41 28 46.425 ;
        RECT 16.65 41 28 46.375 ;
        RECT 16.6 41 28 46.325 ;
        RECT 16.55 41 28 46.275 ;
        RECT 16.45 41 28 46.175 ;
        RECT 16.4 41 28 46.125 ;
        RECT 16.35 41 28 46.075 ;
        RECT 16.3 41 28 46.025 ;
        RECT 16.25 41 28 45.975 ;
        RECT 16.2 41 28 45.925 ;
        RECT 16.15 41 28 45.875 ;
        RECT 16.1 41 28 45.825 ;
        RECT 16.05 41 28 45.775 ;
        RECT 16 41 28 45.725 ;
        RECT 15.95 41 28 45.675 ;
        RECT 15.9 41 28 45.625 ;
        RECT 15.85 41 28 45.575 ;
        RECT 15.8 41 28 45.525 ;
        RECT 15.75 41 28 45.475 ;
        RECT 15.7 41 28 45.425 ;
        RECT 15.65 41 28 45.375 ;
        RECT 15.6 41 28 45.325 ;
        RECT 15.55 41 28 45.275 ;
        RECT 15.5 41 28 45.225 ;
        RECT 15.45 41 28 45.175 ;
        RECT 15.4 41 28 45.125 ;
        RECT 15.35 41 28 45.075 ;
        RECT 15.3 41 28 45.025 ;
        RECT 15.25 41 28 44.975 ;
        RECT 15.2 41 28 44.925 ;
        RECT 15.15 41 28 44.875 ;
        RECT 15.1 41 28 44.825 ;
        RECT 15.05 41 28 44.775 ;
        RECT 15 41 28 44.725 ;
        RECT 14.95 41 28 44.675 ;
        RECT 14.9 41 28 44.625 ;
        RECT 14.85 41 28 44.575 ;
        RECT 14.8 41 28 44.525 ;
        RECT 14.75 41 28 44.475 ;
        RECT 14.7 41 28 44.425 ;
        RECT 14.65 41 28 44.375 ;
        RECT 14.6 41 28 44.325 ;
        RECT 14.55 41 28 44.275 ;
        RECT 14.5 41 28 44.225 ;
        RECT 14.45 41 28 44.175 ;
        RECT 14.4 41 28 44.125 ;
        RECT 14.35 41 28 44.075 ;
        RECT 14.3 41 28 44.025 ;
        RECT 14.25 42.5 33.5 43.975 ;
        RECT 14.2 42.5 33.5 43.925 ;
        RECT 14.15 42.5 33.5 43.875 ;
        RECT 14.1 42.5 33.5 43.825 ;
        RECT 14.05 42.5 33.5 43.775 ;
        RECT 14 42.5 33.5 43.725 ;
        RECT 13.95 42.5 33.5 43.675 ;
        RECT 13.9 42.5 33.5 43.625 ;
        RECT 13.85 42.5 33.5 43.575 ;
        RECT 13.8 42.5 33.5 43.525 ;
        RECT 13.75 42.5 33.5 43.475 ;
        RECT 13.7 42.5 33.5 43.425 ;
        RECT 13.65 42.5 33.5 43.375 ;
        RECT 13.6 42.5 33.5 43.325 ;
        RECT 13.55 42.5 33.5 43.275 ;
        RECT 13.5 42.5 33.5 43.225 ;
        RECT 13.45 42.5 33.5 43.175 ;
        RECT 13.4 42.5 33.5 43.125 ;
        RECT 13.35 42.5 33.5 43.075 ;
        RECT 13.3 42.5 33.5 43.025 ;
        RECT 13.25 42.5 33.5 42.975 ;
        RECT 13.2 42.5 33.5 42.925 ;
        RECT 13.15 42.5 33.5 42.875 ;
        RECT 13.1 42.5 33.5 42.825 ;
        RECT 13.05 42.5 33.5 42.775 ;
        RECT 13 42.5 33.5 42.725 ;
        RECT 12.95 42.5 33.5 42.675 ;
        RECT 12.9 42.5 33.5 42.625 ;
        RECT 12.85 42.5 33.5 42.575 ;
        RECT 4.3 27 12.5 34.025 ;
        RECT 9.5 0 12.5 39.225 ;
        RECT 11.25 34 19.5 40.975 ;
        RECT 11.2 34 19.5 40.925 ;
        RECT 11.15 34 19.5 40.875 ;
        RECT 11.1 34 19.5 40.825 ;
        RECT 11.05 34 19.5 40.775 ;
        RECT 11 34 19.5 40.725 ;
        RECT 10.95 34 19.5 40.675 ;
        RECT 10.9 34 19.5 40.625 ;
        RECT 10.85 34 19.5 40.575 ;
        RECT 10.8 34 19.5 40.525 ;
        RECT 10.75 34 19.5 40.475 ;
        RECT 10.7 34 19.5 40.425 ;
        RECT 10.65 34 19.5 40.375 ;
        RECT 10.6 34 19.5 40.325 ;
        RECT 10.55 34 19.5 40.275 ;
        RECT 10.5 34 19.5 40.225 ;
        RECT 10.45 34 19.5 40.175 ;
        RECT 10.4 34 19.5 40.125 ;
        RECT 10.35 34 19.5 40.075 ;
        RECT 10.3 34 19.5 40.025 ;
        RECT 10.25 34 19.5 39.975 ;
        RECT 10.2 34 19.5 39.925 ;
        RECT 10.15 34 19.5 39.875 ;
        RECT 10.1 34 19.5 39.825 ;
        RECT 10.05 34 19.5 39.775 ;
        RECT 10 34 19.5 39.725 ;
        RECT 9.95 34 19.5 39.675 ;
        RECT 9.9 34 19.5 39.625 ;
        RECT 9.85 34 19.5 39.575 ;
        RECT 9.8 34 19.5 39.525 ;
        RECT 9.75 34 19.5 39.475 ;
        RECT 9.7 34 19.5 39.425 ;
        RECT 9.65 34 19.5 39.375 ;
        RECT 9.6 34 19.5 39.325 ;
        RECT 9.55 34 19.5 39.275 ;
        RECT 9.45 34 19.5 39.175 ;
        RECT 9.4 34 19.5 39.125 ;
        RECT 9.35 34 19.5 39.075 ;
        RECT 9.3 34 19.5 39.025 ;
        RECT 9.25 34 19.5 38.975 ;
        RECT 9.2 34 19.5 38.925 ;
        RECT 9.15 34 19.5 38.875 ;
        RECT 9.1 34 19.5 38.825 ;
        RECT 9.05 34 19.5 38.775 ;
        RECT 9 34 19.5 38.725 ;
        RECT 8.95 34 19.5 38.675 ;
        RECT 8.9 34 19.5 38.625 ;
        RECT 8.85 34 19.5 38.575 ;
        RECT 8.8 34 19.5 38.525 ;
        RECT 8.75 34 19.5 38.475 ;
        RECT 8.7 34 19.5 38.425 ;
        RECT 8.65 34 19.5 38.375 ;
        RECT 8.6 34 19.5 38.325 ;
        RECT 8.55 34 19.5 38.275 ;
        RECT 8.5 34 19.5 38.225 ;
        RECT 8.45 34 19.5 38.175 ;
        RECT 8.4 34 19.5 38.125 ;
        RECT 8.35 34 19.5 38.075 ;
        RECT 8.3 34 19.5 38.025 ;
        RECT 8.25 34 19.5 37.975 ;
        RECT 8.2 34 19.5 37.925 ;
        RECT 8.15 34 19.5 37.875 ;
        RECT 8.1 34 19.5 37.825 ;
        RECT 8.05 34 19.5 37.775 ;
        RECT 8 34 19.5 37.725 ;
        RECT 7.95 34 19.5 37.675 ;
        RECT 7.9 34 19.5 37.625 ;
        RECT 7.85 34 19.5 37.575 ;
        RECT 7.8 34 19.5 37.525 ;
        RECT 7.75 34 19.5 37.475 ;
        RECT 7.7 34 19.5 37.425 ;
        RECT 7.65 34 19.5 37.375 ;
        RECT 7.6 34 19.5 37.325 ;
        RECT 7.55 34 19.5 37.275 ;
        RECT 7.5 34 19.5 37.225 ;
        RECT 7.45 34 19.5 37.175 ;
        RECT 7.4 34 19.5 37.125 ;
        RECT 7.35 34 19.5 37.075 ;
        RECT 7.3 34 19.5 37.025 ;
        RECT 7.25 34 26.5 36.975 ;
        RECT 7.2 34 26.5 36.925 ;
        RECT 7.15 34 26.5 36.875 ;
        RECT 7.1 34 26.5 36.825 ;
        RECT 7.05 34 26.5 36.775 ;
        RECT 7 34 26.5 36.725 ;
        RECT 6.95 34 26.5 36.675 ;
        RECT 6.9 34 26.5 36.625 ;
        RECT 6.85 34 26.5 36.575 ;
        RECT 6.8 34 26.5 36.525 ;
        RECT 6.75 34 26.5 36.475 ;
        RECT 6.7 34 26.5 36.425 ;
        RECT 6.65 34 26.5 36.375 ;
        RECT 6.6 34 26.5 36.325 ;
        RECT 6.55 34 26.5 36.275 ;
        RECT 6.5 34 26.5 36.225 ;
        RECT 6.45 34 26.5 36.175 ;
        RECT 6.4 34 26.5 36.125 ;
        RECT 6.35 34 26.5 36.075 ;
        RECT 6.3 34 26.5 36.025 ;
        RECT 6.25 34 26.5 35.975 ;
        RECT 6.2 34 26.5 35.925 ;
        RECT 6.15 34 26.5 35.875 ;
        RECT 6.1 34 26.5 35.825 ;
        RECT 6.05 34 26.5 35.775 ;
        RECT 6 34 26.5 35.725 ;
        RECT 5.95 34 26.5 35.675 ;
        RECT 5.9 34 26.5 35.625 ;
        RECT 5.85 34 26.5 35.575 ;
        RECT 5.8 34 26.5 35.525 ;
        RECT 5.75 34 26.5 35.475 ;
        RECT 5.7 34 26.5 35.425 ;
        RECT 5.65 34 26.5 35.375 ;
        RECT 5.6 34 26.5 35.325 ;
        RECT 5.55 34 26.5 35.275 ;
        RECT 5.5 34 26.5 35.225 ;
        RECT 1.3 0 5.5 31.025 ;
        RECT 5.45 34 26.5 35.175 ;
        RECT 5.4 34 26.5 35.125 ;
        RECT 5.35 34 26.5 35.075 ;
        RECT 5.3 34 26.5 35.025 ;
        RECT 5.25 34 26.5 34.975 ;
        RECT 5.2 34 26.5 34.925 ;
        RECT 5.15 34 26.5 34.875 ;
        RECT 5.1 34 26.5 34.825 ;
        RECT 5.05 34 26.5 34.775 ;
        RECT 5 34 26.5 34.725 ;
        RECT 4.95 34 26.5 34.675 ;
        RECT 4.9 34 26.5 34.625 ;
        RECT 4.85 34 26.5 34.575 ;
        RECT 4.8 34 26.5 34.525 ;
        RECT 4.75 34 26.5 34.475 ;
        RECT 4.7 34 26.5 34.425 ;
        RECT 4.65 34 26.5 34.375 ;
        RECT 4.6 34 26.5 34.325 ;
        RECT 4.55 34 26.5 34.275 ;
        RECT 4.5 34 26.5 34.225 ;
        RECT 4.45 34 26.5 34.175 ;
        RECT 4.4 34 26.5 34.125 ;
        RECT 4.35 34 26.5 34.075 ;
        RECT 4.25 27 12.5 33.975 ;
        RECT 4.2 27 12.5 33.925 ;
        RECT 4.15 27 12.5 33.875 ;
        RECT 4.1 27 12.5 33.825 ;
        RECT 4.05 27 12.5 33.775 ;
        RECT 4 27 12.5 33.725 ;
        RECT 3.95 27 12.5 33.675 ;
        RECT 3.9 27 12.5 33.625 ;
        RECT 3.85 27 12.5 33.575 ;
        RECT 3.8 27 12.5 33.525 ;
        RECT 3.75 27 12.5 33.475 ;
        RECT 3.7 27 12.5 33.425 ;
        RECT 3.65 27 12.5 33.375 ;
        RECT 3.6 27 12.5 33.325 ;
        RECT 3.55 27 12.5 33.275 ;
        RECT 3.5 27 12.5 33.225 ;
        RECT 3.45 27 12.5 33.175 ;
        RECT 3.4 27 12.5 33.125 ;
        RECT 3.35 27 12.5 33.075 ;
        RECT 3.3 27 12.5 33.025 ;
        RECT 3.25 27 12.5 32.975 ;
        RECT 3.2 27 12.5 32.925 ;
        RECT 3.15 27 12.5 32.875 ;
        RECT 3.1 27 12.5 32.825 ;
        RECT 3.05 27 12.5 32.775 ;
        RECT 3 27 12.5 32.725 ;
        RECT 2.95 27 12.5 32.675 ;
        RECT 2.9 27 12.5 32.625 ;
        RECT 2.85 27 12.5 32.575 ;
        RECT 2.8 27 12.5 32.525 ;
        RECT 2.75 27 12.5 32.475 ;
        RECT 2.7 27 12.5 32.425 ;
        RECT 2.65 27 12.5 32.375 ;
        RECT 2.6 27 12.5 32.325 ;
        RECT 2.55 27 12.5 32.275 ;
        RECT 2.5 27 12.5 32.225 ;
        RECT 2.45 27 12.5 32.175 ;
        RECT 2.4 27 12.5 32.125 ;
        RECT 2.35 27 12.5 32.075 ;
        RECT 2.3 27 12.5 32.025 ;
        RECT 2.25 27 12.5 31.975 ;
        RECT 2.2 27 12.5 31.925 ;
        RECT 2.15 27 12.5 31.875 ;
        RECT 2.1 27 12.5 31.825 ;
        RECT 2.05 27 12.5 31.775 ;
        RECT 2 27 12.5 31.725 ;
        RECT 1.95 27 12.5 31.675 ;
        RECT 1.9 27 12.5 31.625 ;
        RECT 1.85 27 12.5 31.575 ;
        RECT 1.8 27 12.5 31.525 ;
        RECT 1.75 27 12.5 31.475 ;
        RECT 1.7 27 12.5 31.425 ;
        RECT 1.65 27 12.5 31.375 ;
        RECT 1.6 27 12.5 31.325 ;
        RECT 1.55 27 12.5 31.275 ;
        RECT 1.5 27 12.5 31.225 ;
        RECT 1.45 27 12.5 31.175 ;
        RECT 1.4 27 12.5 31.125 ;
        RECT 1.35 27 12.5 31.075 ;
      LAYER M2 ;
        RECT 45 49.5 48 74.7 ;
        RECT 44.95 49.5 48 74.675 ;
        RECT 44.9 49.5 48 74.625 ;
        RECT 44.85 49.5 48 74.575 ;
        RECT 44.8 49.5 48 74.525 ;
        RECT 44.75 49.5 48 74.475 ;
        RECT 44.7 49.5 48 74.425 ;
        RECT 44.65 49.5 48 74.375 ;
        RECT 44.6 49.5 48 74.325 ;
        RECT 44.55 49.5 48 74.275 ;
        RECT 44.5 49.5 48 74.225 ;
        RECT 44.45 62 48 74.175 ;
        RECT 28.3 55 48 58 ;
        RECT 21.3 49.5 48 51 ;
        RECT 44.4 62 48 74.125 ;
        RECT 44.35 62 48 74.075 ;
        RECT 44.3 62 48 74.025 ;
        RECT 44.25 62 48 73.975 ;
        RECT 44.2 62 48 73.925 ;
        RECT 44.15 62 48 73.875 ;
        RECT 44.1 62 48 73.825 ;
        RECT 44.05 62 48 73.775 ;
        RECT 44 62 48 73.725 ;
        RECT 43.95 62 48 73.675 ;
        RECT 43.9 62 48 73.625 ;
        RECT 43.85 62 48 73.575 ;
        RECT 43.8 62 48 73.525 ;
        RECT 43.75 62 48 73.475 ;
        RECT 43.7 62 48 73.425 ;
        RECT 43.65 62 48 73.375 ;
        RECT 43.6 62 48 73.325 ;
        RECT 43.55 62 48 73.275 ;
        RECT 43.5 62 48 73.225 ;
        RECT 43.45 62 48 73.175 ;
        RECT 43.4 62 48 73.125 ;
        RECT 43.35 62 48 73.075 ;
        RECT 43.3 62 48 73.025 ;
        RECT 43.25 62 48 72.975 ;
        RECT 43.2 62 48 72.925 ;
        RECT 43.15 62 48 72.875 ;
        RECT 43.1 62 48 72.825 ;
        RECT 43.05 62 48 72.775 ;
        RECT 43 62 48 72.725 ;
        RECT 42.95 62 48 72.675 ;
        RECT 42.9 62 48 72.625 ;
        RECT 42.85 62 48 72.575 ;
        RECT 42.8 62 48 72.525 ;
        RECT 42.75 62 48 72.475 ;
        RECT 42.7 62 48 72.425 ;
        RECT 42.65 62 48 72.375 ;
        RECT 42.6 62 48 72.325 ;
        RECT 42.55 62 48 72.275 ;
        RECT 42.5 62 48 72.225 ;
        RECT 42.45 62 48 72.175 ;
        RECT 42.4 62 48 72.125 ;
        RECT 42.35 62 48 72.075 ;
        RECT 42.3 62 48 72.025 ;
        RECT 42.25 62 48 71.975 ;
        RECT 42.2 62 48 71.925 ;
        RECT 42.15 62 48 71.875 ;
        RECT 42.1 62 48 71.825 ;
        RECT 42.05 62 48 71.775 ;
        RECT 42 62 48 71.725 ;
        RECT 41.95 62 48 71.675 ;
        RECT 41.9 62 48 71.625 ;
        RECT 41.85 62 48 71.575 ;
        RECT 41.8 62 48 71.525 ;
        RECT 41.75 62 48 71.475 ;
        RECT 41.7 62 48 71.425 ;
        RECT 41.65 62 48 71.375 ;
        RECT 41.6 62 48 71.325 ;
        RECT 41.55 62 48 71.275 ;
        RECT 41.5 62 48 71.225 ;
        RECT 41.45 62 48 71.175 ;
        RECT 41.4 62 48 71.125 ;
        RECT 41.35 62 48 71.075 ;
        RECT 41.3 62 48 71.025 ;
        RECT 41.25 62 48 70.975 ;
        RECT 41.2 62 48 70.925 ;
        RECT 41.15 62 48 70.875 ;
        RECT 41.1 62 48 70.825 ;
        RECT 41.05 62 48 70.775 ;
        RECT 41 62 48 70.725 ;
        RECT 40.95 62 48 70.675 ;
        RECT 40.9 62 48 70.625 ;
        RECT 40.85 62 48 70.575 ;
        RECT 40.8 62 48 70.525 ;
        RECT 40.75 62 48 70.475 ;
        RECT 40.7 62 48 70.425 ;
        RECT 40.65 62 48 70.375 ;
        RECT 40.6 62 48 70.325 ;
        RECT 40.55 62 48 70.275 ;
        RECT 40.5 62 48 70.225 ;
        RECT 32.3 55 40.5 62.025 ;
        RECT 37.5 49.5 40.5 67.225 ;
        RECT 40.45 62 48 70.175 ;
        RECT 40.4 62 48 70.125 ;
        RECT 40.35 62 48 70.075 ;
        RECT 40.3 62 48 70.025 ;
        RECT 40.25 62 48 69.975 ;
        RECT 40.2 62 48 69.925 ;
        RECT 40.15 62 48 69.875 ;
        RECT 40.1 62 48 69.825 ;
        RECT 40.05 62 48 69.775 ;
        RECT 40 62 48 69.725 ;
        RECT 39.95 62 48 69.675 ;
        RECT 39.9 62 48 69.625 ;
        RECT 39.85 62 48 69.575 ;
        RECT 39.8 62 48 69.525 ;
        RECT 39.75 62 48 69.475 ;
        RECT 39.7 62 48 69.425 ;
        RECT 39.65 62 48 69.375 ;
        RECT 39.6 62 48 69.325 ;
        RECT 39.55 62 48 69.275 ;
        RECT 39.5 62 48 69.225 ;
        RECT 39.45 62 48 69.175 ;
        RECT 39.4 62 48 69.125 ;
        RECT 39.35 62 48 69.075 ;
        RECT 39.3 62 48 69.025 ;
        RECT 39.25 62 48 68.975 ;
        RECT 39.2 62 48 68.925 ;
        RECT 39.15 62 48 68.875 ;
        RECT 39.1 62 48 68.825 ;
        RECT 39.05 62 48 68.775 ;
        RECT 39 62 48 68.725 ;
        RECT 38.95 62 48 68.675 ;
        RECT 38.9 62 48 68.625 ;
        RECT 38.85 62 48 68.575 ;
        RECT 38.8 62 48 68.525 ;
        RECT 38.75 62 48 68.475 ;
        RECT 38.7 62 48 68.425 ;
        RECT 38.65 62 48 68.375 ;
        RECT 38.6 62 48 68.325 ;
        RECT 38.55 62 48 68.275 ;
        RECT 38.5 62 48 68.225 ;
        RECT 38.45 62 48 68.175 ;
        RECT 38.4 62 48 68.125 ;
        RECT 38.35 62 48 68.075 ;
        RECT 38.3 62 48 68.025 ;
        RECT 38.25 62 48 67.975 ;
        RECT 38.2 62 48 67.925 ;
        RECT 38.15 62 48 67.875 ;
        RECT 38.1 62 48 67.825 ;
        RECT 38.05 62 48 67.775 ;
        RECT 38 62 48 67.725 ;
        RECT 37.95 62 48 67.675 ;
        RECT 37.9 62 48 67.625 ;
        RECT 37.85 62 48 67.575 ;
        RECT 37.8 62 48 67.525 ;
        RECT 37.75 62 48 67.475 ;
        RECT 37.7 62 48 67.425 ;
        RECT 37.65 62 48 67.375 ;
        RECT 37.6 62 48 67.325 ;
        RECT 37.55 62 48 67.275 ;
        RECT 37.45 62 48 67.175 ;
        RECT 37.4 62 48 67.125 ;
        RECT 37.35 62 48 67.075 ;
        RECT 37.3 62 48 67.025 ;
        RECT 37.25 62 48 66.975 ;
        RECT 37.2 62 48 66.925 ;
        RECT 37.15 62 48 66.875 ;
        RECT 37.1 62 48 66.825 ;
        RECT 37.05 62 48 66.775 ;
        RECT 37 62 48 66.725 ;
        RECT 19.8 49.475 37 49.525 ;
        RECT 36.95 62 48 66.675 ;
        RECT 19.75 49.425 36.95 49.475 ;
        RECT 36.9 62 48 66.625 ;
        RECT 19.7 49.375 36.9 49.425 ;
        RECT 36.85 62 48 66.575 ;
        RECT 19.65 49.325 36.85 49.375 ;
        RECT 36.8 62 48 66.525 ;
        RECT 19.6 49.275 36.8 49.325 ;
        RECT 36.75 62 48 66.475 ;
        RECT 19.55 49.225 36.75 49.275 ;
        RECT 36.7 62 48 66.425 ;
        RECT 19.5 49.175 36.7 49.225 ;
        RECT 36.65 62 48 66.375 ;
        RECT 19.45 49.125 36.65 49.175 ;
        RECT 36.6 62 48 66.325 ;
        RECT 19.4 49.075 36.6 49.125 ;
        RECT 36.55 62 48 66.275 ;
        RECT 19.35 49.025 36.55 49.075 ;
        RECT 36.5 62 48 66.225 ;
        RECT 19.3 48.975 36.5 49.025 ;
        RECT 36.45 62 48 66.175 ;
        RECT 19.25 48.925 36.45 48.975 ;
        RECT 36.4 62 48 66.125 ;
        RECT 19.2 48.875 36.4 48.925 ;
        RECT 36.35 62 48 66.075 ;
        RECT 19.15 48.825 36.35 48.875 ;
        RECT 36.3 62 48 66.025 ;
        RECT 19.1 48.775 36.3 48.825 ;
        RECT 36.25 62 48 65.975 ;
        RECT 19.05 48.725 36.25 48.775 ;
        RECT 36.2 62 48 65.925 ;
        RECT 19 48.675 36.2 48.725 ;
        RECT 36.15 62 48 65.875 ;
        RECT 18.95 48.625 36.15 48.675 ;
        RECT 36.1 62 48 65.825 ;
        RECT 18.9 48.575 36.1 48.625 ;
        RECT 36.05 62 48 65.775 ;
        RECT 18.85 48.525 36.05 48.575 ;
        RECT 36 62 48 65.725 ;
        RECT 18.8 48.475 36 48.525 ;
        RECT 35.95 62 48 65.675 ;
        RECT 18.75 48.425 35.95 48.475 ;
        RECT 35.9 62 48 65.625 ;
        RECT 18.7 48.375 35.9 48.425 ;
        RECT 35.85 62 48 65.575 ;
        RECT 18.65 48.325 35.85 48.375 ;
        RECT 35.8 62 48 65.525 ;
        RECT 18.6 48.275 35.8 48.325 ;
        RECT 35.75 62 48 65.475 ;
        RECT 18.55 48.225 35.75 48.275 ;
        RECT 35.7 62 48 65.425 ;
        RECT 18.5 48.175 35.7 48.225 ;
        RECT 35.65 62 48 65.375 ;
        RECT 18.45 48.125 35.65 48.175 ;
        RECT 35.6 62 48 65.325 ;
        RECT 18.4 48.075 35.6 48.125 ;
        RECT 35.55 62 48 65.275 ;
        RECT 18.35 48.025 35.55 48.075 ;
        RECT 35.5 62 48 65.225 ;
        RECT 32 47.975 35.5 51 ;
        RECT 35.45 62 48 65.175 ;
        RECT 32 47.925 35.45 51 ;
        RECT 35.4 62 48 65.125 ;
        RECT 32 47.875 35.4 51 ;
        RECT 35.35 62 48 65.075 ;
        RECT 32 47.825 35.35 51 ;
        RECT 35.3 62 48 65.025 ;
        RECT 32 47.775 35.3 51 ;
        RECT 35.25 62 48 64.975 ;
        RECT 32 47.725 35.25 51 ;
        RECT 35.2 62 48 64.925 ;
        RECT 32 47.675 35.2 51 ;
        RECT 35.15 62 48 64.875 ;
        RECT 32 47.625 35.15 51 ;
        RECT 35.1 62 48 64.825 ;
        RECT 32 47.575 35.1 51 ;
        RECT 35.05 62 48 64.775 ;
        RECT 32 47.525 35.05 51 ;
        RECT 35 62 48 64.725 ;
        RECT 32 47.475 35 51 ;
        RECT 34.95 62 48 64.675 ;
        RECT 32 47.425 34.95 51 ;
        RECT 34.9 62 48 64.625 ;
        RECT 32 47.375 34.9 51 ;
        RECT 34.85 62 48 64.575 ;
        RECT 32 47.325 34.85 51 ;
        RECT 34.8 62 48 64.525 ;
        RECT 32 47.275 34.8 51 ;
        RECT 34.75 62 48 64.475 ;
        RECT 32 47.225 34.75 51 ;
        RECT 34.7 62 48 64.425 ;
        RECT 32 47.175 34.7 51 ;
        RECT 34.65 62 48 64.375 ;
        RECT 32 47.125 34.65 51 ;
        RECT 34.6 62 48 64.325 ;
        RECT 32 47.075 34.6 51 ;
        RECT 34.55 62 48 64.275 ;
        RECT 32 47.025 34.55 51 ;
        RECT 34.5 62 48 64.225 ;
        RECT 32 46.975 34.5 51 ;
        RECT 34.45 62 48 64.175 ;
        RECT 32 46.925 34.45 51 ;
        RECT 34.4 62 48 64.125 ;
        RECT 32 46.875 34.4 51 ;
        RECT 34.35 62 48 64.075 ;
        RECT 32 46.825 34.35 51 ;
        RECT 34.3 62 48 64.025 ;
        RECT 32 46.775 34.3 51 ;
        RECT 34.25 62 48 63.975 ;
        RECT 32 46.725 34.25 51 ;
        RECT 34.2 62 48 63.925 ;
        RECT 32 46.675 34.2 51 ;
        RECT 34.15 62 48 63.875 ;
        RECT 32 46.625 34.15 51 ;
        RECT 34.1 62 48 63.825 ;
        RECT 32 46.575 34.1 51 ;
        RECT 34.05 62 48 63.775 ;
        RECT 32 46.525 34.05 51 ;
        RECT 34 62 48 63.725 ;
        RECT 32 46.475 34 51 ;
        RECT 33.95 62 48 63.675 ;
        RECT 32 46.425 33.95 51 ;
        RECT 33.9 62 48 63.625 ;
        RECT 32 46.375 33.9 51 ;
        RECT 33.85 62 48 63.575 ;
        RECT 32 46.325 33.85 51 ;
        RECT 33.8 62 48 63.525 ;
        RECT 32 46.275 33.8 51 ;
        RECT 33.75 62 48 63.475 ;
        RECT 32 46.225 33.75 51 ;
        RECT 33.7 62 48 63.425 ;
        RECT 32 46.175 33.7 51 ;
        RECT 33.65 62 48 63.375 ;
        RECT 32 46.125 33.65 51 ;
        RECT 33.6 62 48 63.325 ;
        RECT 32 46.075 33.6 51 ;
        RECT 33.55 62 48 63.275 ;
        RECT 32 46.025 33.55 51 ;
        RECT 33.5 62 48 63.225 ;
        RECT 25.3 48 33.5 55.025 ;
        RECT 32 42.5 33.5 61.725 ;
        RECT 33.45 62 48 63.175 ;
        RECT 33.4 62 48 63.125 ;
        RECT 33.35 62 48 63.075 ;
        RECT 33.3 62 48 63.025 ;
        RECT 33.25 62 48 62.975 ;
        RECT 33.2 62 48 62.925 ;
        RECT 33.15 62 48 62.875 ;
        RECT 33.1 62 48 62.825 ;
        RECT 33.05 62 48 62.775 ;
        RECT 33 62 48 62.725 ;
        RECT 32.95 62 48 62.675 ;
        RECT 32.9 62 48 62.625 ;
        RECT 32.85 62 48 62.575 ;
        RECT 32.8 62 48 62.525 ;
        RECT 32.75 62 48 62.475 ;
        RECT 32.7 62 48 62.425 ;
        RECT 32.65 62 48 62.375 ;
        RECT 32.6 62 48 62.325 ;
        RECT 32.55 62 48 62.275 ;
        RECT 32.5 62 48 62.225 ;
        RECT 32.45 62 48 62.175 ;
        RECT 32.4 62 48 62.125 ;
        RECT 32.35 62 48 62.075 ;
        RECT 32.25 55 40.5 61.975 ;
        RECT 32.2 55 40.5 61.925 ;
        RECT 32.15 55 40.5 61.875 ;
        RECT 32.1 55 40.5 61.825 ;
        RECT 32.05 55 40.5 61.775 ;
        RECT 31.95 55 40.5 61.675 ;
        RECT 14.3 42.5 33.5 44 ;
        RECT 31.9 55 40.5 61.625 ;
        RECT 31.85 55 40.5 61.575 ;
        RECT 31.8 55 40.5 61.525 ;
        RECT 31.75 55 40.5 61.475 ;
        RECT 31.7 55 40.5 61.425 ;
        RECT 31.65 55 40.5 61.375 ;
        RECT 31.6 55 40.5 61.325 ;
        RECT 31.55 55 40.5 61.275 ;
        RECT 31.5 55 40.5 61.225 ;
        RECT 31.45 55 40.5 61.175 ;
        RECT 31.4 55 40.5 61.125 ;
        RECT 31.35 55 40.5 61.075 ;
        RECT 31.3 55 40.5 61.025 ;
        RECT 31.25 55 40.5 60.975 ;
        RECT 31.2 55 40.5 60.925 ;
        RECT 31.15 55 40.5 60.875 ;
        RECT 31.1 55 40.5 60.825 ;
        RECT 31.05 55 40.5 60.775 ;
        RECT 31 55 40.5 60.725 ;
        RECT 30.95 55 40.5 60.675 ;
        RECT 30.9 55 40.5 60.625 ;
        RECT 30.85 55 40.5 60.575 ;
        RECT 30.8 55 40.5 60.525 ;
        RECT 30.75 55 40.5 60.475 ;
        RECT 30.7 55 40.5 60.425 ;
        RECT 30.65 55 40.5 60.375 ;
        RECT 30.6 55 40.5 60.325 ;
        RECT 30.55 55 40.5 60.275 ;
        RECT 30.5 55 40.5 60.225 ;
        RECT 30.45 55 40.5 60.175 ;
        RECT 30.4 55 40.5 60.125 ;
        RECT 30.35 55 40.5 60.075 ;
        RECT 30.3 55 40.5 60.025 ;
        RECT 30.25 55 40.5 59.975 ;
        RECT 30.2 55 40.5 59.925 ;
        RECT 30.15 55 40.5 59.875 ;
        RECT 30.1 55 40.5 59.825 ;
        RECT 30.05 55 40.5 59.775 ;
        RECT 30 55 40.5 59.725 ;
        RECT 12.8 42.475 30 42.525 ;
        RECT 29.95 55 40.5 59.675 ;
        RECT 12.75 42.425 29.95 42.475 ;
        RECT 29.9 55 40.5 59.625 ;
        RECT 12.7 42.375 29.9 42.425 ;
        RECT 29.85 55 40.5 59.575 ;
        RECT 12.65 42.325 29.85 42.375 ;
        RECT 29.8 55 40.5 59.525 ;
        RECT 12.6 42.275 29.8 42.325 ;
        RECT 29.75 55 40.5 59.475 ;
        RECT 12.55 42.225 29.75 42.275 ;
        RECT 29.7 55 40.5 59.425 ;
        RECT 12.5 42.175 29.7 42.225 ;
        RECT 29.65 55 40.5 59.375 ;
        RECT 12.45 42.125 29.65 42.175 ;
        RECT 29.6 55 40.5 59.325 ;
        RECT 12.4 42.075 29.6 42.125 ;
        RECT 29.55 55 40.5 59.275 ;
        RECT 12.35 42.025 29.55 42.075 ;
        RECT 29.5 55 40.5 59.225 ;
        RECT 12.3 41.975 29.5 42.025 ;
        RECT 29.45 55 40.5 59.175 ;
        RECT 12.25 41.925 29.45 41.975 ;
        RECT 29.4 55 40.5 59.125 ;
        RECT 12.2 41.875 29.4 41.925 ;
        RECT 29.35 55 40.5 59.075 ;
        RECT 12.15 41.825 29.35 41.875 ;
        RECT 29.3 55 40.5 59.025 ;
        RECT 12.1 41.775 29.3 41.825 ;
        RECT 29.25 55 40.5 58.975 ;
        RECT 12.05 41.725 29.25 41.775 ;
        RECT 29.2 55 40.5 58.925 ;
        RECT 12 41.675 29.2 41.725 ;
        RECT 29.15 55 40.5 58.875 ;
        RECT 11.95 41.625 29.15 41.675 ;
        RECT 29.1 55 40.5 58.825 ;
        RECT 11.9 41.575 29.1 41.625 ;
        RECT 29.05 55 40.5 58.775 ;
        RECT 11.85 41.525 29.05 41.575 ;
        RECT 29 55 40.5 58.725 ;
        RECT 11.8 41.475 29 41.525 ;
        RECT 28.95 55 40.5 58.675 ;
        RECT 11.75 41.425 28.95 41.475 ;
        RECT 28.9 55 40.5 58.625 ;
        RECT 11.7 41.375 28.9 41.425 ;
        RECT 28.85 55 40.5 58.575 ;
        RECT 11.65 41.325 28.85 41.375 ;
        RECT 28.8 55 40.5 58.525 ;
        RECT 11.6 41.275 28.8 41.325 ;
        RECT 28.75 55 40.5 58.475 ;
        RECT 11.55 41.225 28.75 41.275 ;
        RECT 28.7 55 40.5 58.425 ;
        RECT 11.5 41.175 28.7 41.225 ;
        RECT 28.65 55 40.5 58.375 ;
        RECT 11.45 41.125 28.65 41.175 ;
        RECT 28.6 55 40.5 58.325 ;
        RECT 11.4 41.075 28.6 41.125 ;
        RECT 28.55 55 40.5 58.275 ;
        RECT 11.35 41.025 28.55 41.075 ;
        RECT 28.5 55 40.5 58.225 ;
        RECT 23.5 40.975 28.5 44 ;
        RECT 28.45 55 40.5 58.175 ;
        RECT 23.5 40.925 28.45 44 ;
        RECT 28.4 55 40.5 58.125 ;
        RECT 23.5 40.875 28.4 44 ;
        RECT 28.35 55 40.5 58.075 ;
        RECT 23.5 40.825 28.35 44 ;
        RECT 28.3 55 40.5 58.025 ;
        RECT 23.5 40.775 28.3 44 ;
        RECT 28.25 55 48 57.975 ;
        RECT 23.5 40.725 28.25 44 ;
        RECT 28.2 55 48 57.925 ;
        RECT 23.5 40.675 28.2 44 ;
        RECT 28.15 55 48 57.875 ;
        RECT 23.5 40.625 28.15 44 ;
        RECT 28.1 55 48 57.825 ;
        RECT 23.5 40.575 28.1 44 ;
        RECT 28.05 55 48 57.775 ;
        RECT 23.5 40.525 28.05 44 ;
        RECT 28 55 48 57.725 ;
        RECT 18.3 41 28 48.025 ;
        RECT 23.5 40.475 28 53.225 ;
        RECT 27.95 55 48 57.675 ;
        RECT 23.5 40.425 27.95 53.225 ;
        RECT 27.9 55 48 57.625 ;
        RECT 23.5 40.375 27.9 53.225 ;
        RECT 27.85 55 48 57.575 ;
        RECT 23.5 40.325 27.85 53.225 ;
        RECT 27.8 55 48 57.525 ;
        RECT 23.5 40.275 27.8 53.225 ;
        RECT 27.75 55 48 57.475 ;
        RECT 23.5 40.225 27.75 53.225 ;
        RECT 27.7 55 48 57.425 ;
        RECT 23.5 40.175 27.7 53.225 ;
        RECT 27.65 55 48 57.375 ;
        RECT 23.5 40.125 27.65 53.225 ;
        RECT 27.6 55 48 57.325 ;
        RECT 23.5 40.075 27.6 53.225 ;
        RECT 27.55 55 48 57.275 ;
        RECT 23.5 40.025 27.55 53.225 ;
        RECT 27.5 55 48 57.225 ;
        RECT 23.5 39.975 27.5 53.225 ;
        RECT 27.45 55 48 57.175 ;
        RECT 23.5 39.925 27.45 53.225 ;
        RECT 27.4 55 48 57.125 ;
        RECT 23.5 39.875 27.4 53.225 ;
        RECT 27.35 55 48 57.075 ;
        RECT 23.5 39.825 27.35 53.225 ;
        RECT 27.3 55 48 57.025 ;
        RECT 23.5 39.775 27.3 53.225 ;
        RECT 27.25 55 48 56.975 ;
        RECT 23.5 39.725 27.25 53.225 ;
        RECT 27.2 55 48 56.925 ;
        RECT 23.5 39.675 27.2 53.225 ;
        RECT 27.15 55 48 56.875 ;
        RECT 23.5 39.625 27.15 53.225 ;
        RECT 27.1 55 48 56.825 ;
        RECT 23.5 39.575 27.1 53.225 ;
        RECT 27.05 55 48 56.775 ;
        RECT 23.5 39.525 27.05 53.225 ;
        RECT 27 55 48 56.725 ;
        RECT 23.5 39.475 27 53.225 ;
        RECT 26.95 55 48 56.675 ;
        RECT 23.5 39.425 26.95 53.225 ;
        RECT 26.9 55 48 56.625 ;
        RECT 23.5 39.375 26.9 53.225 ;
        RECT 26.85 55 48 56.575 ;
        RECT 23.5 39.325 26.85 53.225 ;
        RECT 26.8 55 48 56.525 ;
        RECT 23.5 39.275 26.8 53.225 ;
        RECT 26.75 55 48 56.475 ;
        RECT 23.5 39.225 26.75 53.225 ;
        RECT 26.7 55 48 56.425 ;
        RECT 23.5 39.175 26.7 53.225 ;
        RECT 26.65 55 48 56.375 ;
        RECT 23.5 39.125 26.65 53.225 ;
        RECT 26.6 55 48 56.325 ;
        RECT 23.5 39.075 26.6 53.225 ;
        RECT 26.55 55 48 56.275 ;
        RECT 23.5 39.025 26.55 53.225 ;
        RECT 26.5 55 48 56.225 ;
        RECT 23.5 0 26.5 53.225 ;
        RECT 26.45 55 48 56.175 ;
        RECT 26.4 55 48 56.125 ;
        RECT 26.35 55 48 56.075 ;
        RECT 26.3 55 48 56.025 ;
        RECT 26.25 55 48 55.975 ;
        RECT 26.2 55 48 55.925 ;
        RECT 26.15 55 48 55.875 ;
        RECT 26.1 55 48 55.825 ;
        RECT 26.05 55 48 55.775 ;
        RECT 26 55 48 55.725 ;
        RECT 25.95 55 48 55.675 ;
        RECT 25.9 55 48 55.625 ;
        RECT 25.85 55 48 55.575 ;
        RECT 25.8 55 48 55.525 ;
        RECT 25.75 55 48 55.475 ;
        RECT 25.7 55 48 55.425 ;
        RECT 25.65 55 48 55.375 ;
        RECT 25.6 55 48 55.325 ;
        RECT 25.55 55 48 55.275 ;
        RECT 25.5 55 48 55.225 ;
        RECT 25.45 55 48 55.175 ;
        RECT 25.4 55 48 55.125 ;
        RECT 25.35 55 48 55.075 ;
        RECT 25.25 48 33.5 54.975 ;
        RECT 25.2 48 33.5 54.925 ;
        RECT 25.15 48 33.5 54.875 ;
        RECT 25.1 48 33.5 54.825 ;
        RECT 25.05 48 33.5 54.775 ;
        RECT 25 48 33.5 54.725 ;
        RECT 24.95 48 33.5 54.675 ;
        RECT 24.9 48 33.5 54.625 ;
        RECT 24.85 48 33.5 54.575 ;
        RECT 24.8 48 33.5 54.525 ;
        RECT 24.75 48 33.5 54.475 ;
        RECT 24.7 48 33.5 54.425 ;
        RECT 24.65 48 33.5 54.375 ;
        RECT 24.6 48 33.5 54.325 ;
        RECT 24.55 48 33.5 54.275 ;
        RECT 24.5 48 33.5 54.225 ;
        RECT 24.45 48 33.5 54.175 ;
        RECT 24.4 48 33.5 54.125 ;
        RECT 24.35 48 33.5 54.075 ;
        RECT 24.3 48 33.5 54.025 ;
        RECT 24.25 48 33.5 53.975 ;
        RECT 24.2 48 33.5 53.925 ;
        RECT 24.15 48 33.5 53.875 ;
        RECT 24.1 48 33.5 53.825 ;
        RECT 24.05 48 33.5 53.775 ;
        RECT 24 48 33.5 53.725 ;
        RECT 23.95 48 33.5 53.675 ;
        RECT 23.9 48 33.5 53.625 ;
        RECT 23.85 48 33.5 53.575 ;
        RECT 23.8 48 33.5 53.525 ;
        RECT 23.75 48 33.5 53.475 ;
        RECT 23.7 48 33.5 53.425 ;
        RECT 23.65 48 33.5 53.375 ;
        RECT 23.6 48 33.5 53.325 ;
        RECT 23.55 48 33.5 53.275 ;
        RECT 23.45 48 33.5 53.175 ;
        RECT 7.3 34 26.5 37 ;
        RECT 1.3 27 26.5 30 ;
        RECT 1.3 20 26.5 23 ;
        RECT 1.3 13 26.5 16 ;
        RECT 1.3 6 26.5 9 ;
        RECT 1.3 0 26.5 2 ;
        RECT 23.4 48 33.5 53.125 ;
        RECT 23.35 48 33.5 53.075 ;
        RECT 23.3 48 33.5 53.025 ;
        RECT 23.25 48 33.5 52.975 ;
        RECT 23.2 48 33.5 52.925 ;
        RECT 23.15 48 33.5 52.875 ;
        RECT 23.1 48 33.5 52.825 ;
        RECT 23.05 48 33.5 52.775 ;
        RECT 23 48 33.5 52.725 ;
        RECT 22.95 48 33.5 52.675 ;
        RECT 22.9 48 33.5 52.625 ;
        RECT 22.85 48 33.5 52.575 ;
        RECT 22.8 48 33.5 52.525 ;
        RECT 22.75 48 33.5 52.475 ;
        RECT 22.7 48 33.5 52.425 ;
        RECT 22.65 48 33.5 52.375 ;
        RECT 22.6 48 33.5 52.325 ;
        RECT 22.55 48 33.5 52.275 ;
        RECT 22.5 48 33.5 52.225 ;
        RECT 22.45 48 33.5 52.175 ;
        RECT 22.4 48 33.5 52.125 ;
        RECT 22.35 48 33.5 52.075 ;
        RECT 22.3 48 33.5 52.025 ;
        RECT 22.25 48 33.5 51.975 ;
        RECT 22.2 48 33.5 51.925 ;
        RECT 22.15 48 33.5 51.875 ;
        RECT 22.1 48 33.5 51.825 ;
        RECT 22.05 48 33.5 51.775 ;
        RECT 22 48 33.5 51.725 ;
        RECT 21.95 48 33.5 51.675 ;
        RECT 21.9 48 33.5 51.625 ;
        RECT 21.85 48 33.5 51.575 ;
        RECT 21.8 48 33.5 51.525 ;
        RECT 21.75 48 33.5 51.475 ;
        RECT 21.7 48 33.5 51.425 ;
        RECT 21.65 48 33.5 51.375 ;
        RECT 21.6 48 33.5 51.325 ;
        RECT 21.55 48 33.5 51.275 ;
        RECT 21.5 48 33.5 51.225 ;
        RECT 21.45 48 33.5 51.175 ;
        RECT 21.4 48 33.5 51.125 ;
        RECT 21.35 48 33.5 51.075 ;
        RECT 21.3 48 33.5 51.025 ;
        RECT 21.25 49.5 48 50.975 ;
        RECT 21.2 49.5 48 50.925 ;
        RECT 21.15 49.5 48 50.875 ;
        RECT 21.1 49.5 48 50.825 ;
        RECT 21.05 49.5 48 50.775 ;
        RECT 21 49.5 48 50.725 ;
        RECT 20.95 49.5 48 50.675 ;
        RECT 20.9 49.5 48 50.625 ;
        RECT 20.85 49.5 48 50.575 ;
        RECT 20.8 49.5 48 50.525 ;
        RECT 20.75 49.5 48 50.475 ;
        RECT 20.7 49.5 48 50.425 ;
        RECT 20.65 49.5 48 50.375 ;
        RECT 20.6 49.5 48 50.325 ;
        RECT 20.55 49.5 48 50.275 ;
        RECT 20.5 49.5 48 50.225 ;
        RECT 20.45 49.5 48 50.175 ;
        RECT 20.4 49.5 48 50.125 ;
        RECT 20.35 49.5 48 50.075 ;
        RECT 20.3 49.5 48 50.025 ;
        RECT 20.25 49.5 48 49.975 ;
        RECT 20.2 49.5 48 49.925 ;
        RECT 20.15 49.5 48 49.875 ;
        RECT 20.1 49.5 48 49.825 ;
        RECT 20.05 49.5 48 49.775 ;
        RECT 20 49.5 48 49.725 ;
        RECT 19.95 49.5 48 49.675 ;
        RECT 19.9 49.5 48 49.625 ;
        RECT 19.85 49.5 48 49.575 ;
        RECT 11.3 34 19.5 41.025 ;
        RECT 16.5 0 19.5 46.225 ;
        RECT 18.25 41 28 47.975 ;
        RECT 18.2 41 28 47.925 ;
        RECT 18.15 41 28 47.875 ;
        RECT 18.1 41 28 47.825 ;
        RECT 18.05 41 28 47.775 ;
        RECT 18 41 28 47.725 ;
        RECT 17.95 41 28 47.675 ;
        RECT 17.9 41 28 47.625 ;
        RECT 17.85 41 28 47.575 ;
        RECT 17.8 41 28 47.525 ;
        RECT 17.75 41 28 47.475 ;
        RECT 17.7 41 28 47.425 ;
        RECT 17.65 41 28 47.375 ;
        RECT 17.6 41 28 47.325 ;
        RECT 17.55 41 28 47.275 ;
        RECT 17.5 41 28 47.225 ;
        RECT 17.45 41 28 47.175 ;
        RECT 17.4 41 28 47.125 ;
        RECT 17.35 41 28 47.075 ;
        RECT 17.3 41 28 47.025 ;
        RECT 17.25 41 28 46.975 ;
        RECT 17.2 41 28 46.925 ;
        RECT 17.15 41 28 46.875 ;
        RECT 17.1 41 28 46.825 ;
        RECT 17.05 41 28 46.775 ;
        RECT 17 41 28 46.725 ;
        RECT 16.95 41 28 46.675 ;
        RECT 16.9 41 28 46.625 ;
        RECT 16.85 41 28 46.575 ;
        RECT 16.8 41 28 46.525 ;
        RECT 16.75 41 28 46.475 ;
        RECT 16.7 41 28 46.425 ;
        RECT 16.65 41 28 46.375 ;
        RECT 16.6 41 28 46.325 ;
        RECT 16.55 41 28 46.275 ;
        RECT 16.45 41 28 46.175 ;
        RECT 16.4 41 28 46.125 ;
        RECT 16.35 41 28 46.075 ;
        RECT 16.3 41 28 46.025 ;
        RECT 16.25 41 28 45.975 ;
        RECT 16.2 41 28 45.925 ;
        RECT 16.15 41 28 45.875 ;
        RECT 16.1 41 28 45.825 ;
        RECT 16.05 41 28 45.775 ;
        RECT 16 41 28 45.725 ;
        RECT 15.95 41 28 45.675 ;
        RECT 15.9 41 28 45.625 ;
        RECT 15.85 41 28 45.575 ;
        RECT 15.8 41 28 45.525 ;
        RECT 15.75 41 28 45.475 ;
        RECT 15.7 41 28 45.425 ;
        RECT 15.65 41 28 45.375 ;
        RECT 15.6 41 28 45.325 ;
        RECT 15.55 41 28 45.275 ;
        RECT 15.5 41 28 45.225 ;
        RECT 15.45 41 28 45.175 ;
        RECT 15.4 41 28 45.125 ;
        RECT 15.35 41 28 45.075 ;
        RECT 15.3 41 28 45.025 ;
        RECT 15.25 41 28 44.975 ;
        RECT 15.2 41 28 44.925 ;
        RECT 15.15 41 28 44.875 ;
        RECT 15.1 41 28 44.825 ;
        RECT 15.05 41 28 44.775 ;
        RECT 15 41 28 44.725 ;
        RECT 14.95 41 28 44.675 ;
        RECT 14.9 41 28 44.625 ;
        RECT 14.85 41 28 44.575 ;
        RECT 14.8 41 28 44.525 ;
        RECT 14.75 41 28 44.475 ;
        RECT 14.7 41 28 44.425 ;
        RECT 14.65 41 28 44.375 ;
        RECT 14.6 41 28 44.325 ;
        RECT 14.55 41 28 44.275 ;
        RECT 14.5 41 28 44.225 ;
        RECT 14.45 41 28 44.175 ;
        RECT 14.4 41 28 44.125 ;
        RECT 14.35 41 28 44.075 ;
        RECT 14.3 41 28 44.025 ;
        RECT 14.25 42.5 33.5 43.975 ;
        RECT 14.2 42.5 33.5 43.925 ;
        RECT 14.15 42.5 33.5 43.875 ;
        RECT 14.1 42.5 33.5 43.825 ;
        RECT 14.05 42.5 33.5 43.775 ;
        RECT 14 42.5 33.5 43.725 ;
        RECT 13.95 42.5 33.5 43.675 ;
        RECT 13.9 42.5 33.5 43.625 ;
        RECT 13.85 42.5 33.5 43.575 ;
        RECT 13.8 42.5 33.5 43.525 ;
        RECT 13.75 42.5 33.5 43.475 ;
        RECT 13.7 42.5 33.5 43.425 ;
        RECT 13.65 42.5 33.5 43.375 ;
        RECT 13.6 42.5 33.5 43.325 ;
        RECT 13.55 42.5 33.5 43.275 ;
        RECT 13.5 42.5 33.5 43.225 ;
        RECT 13.45 42.5 33.5 43.175 ;
        RECT 13.4 42.5 33.5 43.125 ;
        RECT 13.35 42.5 33.5 43.075 ;
        RECT 13.3 42.5 33.5 43.025 ;
        RECT 13.25 42.5 33.5 42.975 ;
        RECT 13.2 42.5 33.5 42.925 ;
        RECT 13.15 42.5 33.5 42.875 ;
        RECT 13.1 42.5 33.5 42.825 ;
        RECT 13.05 42.5 33.5 42.775 ;
        RECT 13 42.5 33.5 42.725 ;
        RECT 12.95 42.5 33.5 42.675 ;
        RECT 12.9 42.5 33.5 42.625 ;
        RECT 12.85 42.5 33.5 42.575 ;
        RECT 4.3 27 12.5 34.025 ;
        RECT 9.5 0 12.5 39.225 ;
        RECT 11.25 34 19.5 40.975 ;
        RECT 11.2 34 19.5 40.925 ;
        RECT 11.15 34 19.5 40.875 ;
        RECT 11.1 34 19.5 40.825 ;
        RECT 11.05 34 19.5 40.775 ;
        RECT 11 34 19.5 40.725 ;
        RECT 10.95 34 19.5 40.675 ;
        RECT 10.9 34 19.5 40.625 ;
        RECT 10.85 34 19.5 40.575 ;
        RECT 10.8 34 19.5 40.525 ;
        RECT 10.75 34 19.5 40.475 ;
        RECT 10.7 34 19.5 40.425 ;
        RECT 10.65 34 19.5 40.375 ;
        RECT 10.6 34 19.5 40.325 ;
        RECT 10.55 34 19.5 40.275 ;
        RECT 10.5 34 19.5 40.225 ;
        RECT 10.45 34 19.5 40.175 ;
        RECT 10.4 34 19.5 40.125 ;
        RECT 10.35 34 19.5 40.075 ;
        RECT 10.3 34 19.5 40.025 ;
        RECT 10.25 34 19.5 39.975 ;
        RECT 10.2 34 19.5 39.925 ;
        RECT 10.15 34 19.5 39.875 ;
        RECT 10.1 34 19.5 39.825 ;
        RECT 10.05 34 19.5 39.775 ;
        RECT 10 34 19.5 39.725 ;
        RECT 9.95 34 19.5 39.675 ;
        RECT 9.9 34 19.5 39.625 ;
        RECT 9.85 34 19.5 39.575 ;
        RECT 9.8 34 19.5 39.525 ;
        RECT 9.75 34 19.5 39.475 ;
        RECT 9.7 34 19.5 39.425 ;
        RECT 9.65 34 19.5 39.375 ;
        RECT 9.6 34 19.5 39.325 ;
        RECT 9.55 34 19.5 39.275 ;
        RECT 9.45 34 19.5 39.175 ;
        RECT 9.4 34 19.5 39.125 ;
        RECT 9.35 34 19.5 39.075 ;
        RECT 9.3 34 19.5 39.025 ;
        RECT 9.25 34 19.5 38.975 ;
        RECT 9.2 34 19.5 38.925 ;
        RECT 9.15 34 19.5 38.875 ;
        RECT 9.1 34 19.5 38.825 ;
        RECT 9.05 34 19.5 38.775 ;
        RECT 9 34 19.5 38.725 ;
        RECT 8.95 34 19.5 38.675 ;
        RECT 8.9 34 19.5 38.625 ;
        RECT 8.85 34 19.5 38.575 ;
        RECT 8.8 34 19.5 38.525 ;
        RECT 8.75 34 19.5 38.475 ;
        RECT 8.7 34 19.5 38.425 ;
        RECT 8.65 34 19.5 38.375 ;
        RECT 8.6 34 19.5 38.325 ;
        RECT 8.55 34 19.5 38.275 ;
        RECT 8.5 34 19.5 38.225 ;
        RECT 8.45 34 19.5 38.175 ;
        RECT 8.4 34 19.5 38.125 ;
        RECT 8.35 34 19.5 38.075 ;
        RECT 8.3 34 19.5 38.025 ;
        RECT 8.25 34 19.5 37.975 ;
        RECT 8.2 34 19.5 37.925 ;
        RECT 8.15 34 19.5 37.875 ;
        RECT 8.1 34 19.5 37.825 ;
        RECT 8.05 34 19.5 37.775 ;
        RECT 8 34 19.5 37.725 ;
        RECT 7.95 34 19.5 37.675 ;
        RECT 7.9 34 19.5 37.625 ;
        RECT 7.85 34 19.5 37.575 ;
        RECT 7.8 34 19.5 37.525 ;
        RECT 7.75 34 19.5 37.475 ;
        RECT 7.7 34 19.5 37.425 ;
        RECT 7.65 34 19.5 37.375 ;
        RECT 7.6 34 19.5 37.325 ;
        RECT 7.55 34 19.5 37.275 ;
        RECT 7.5 34 19.5 37.225 ;
        RECT 7.45 34 19.5 37.175 ;
        RECT 7.4 34 19.5 37.125 ;
        RECT 7.35 34 19.5 37.075 ;
        RECT 7.3 34 19.5 37.025 ;
        RECT 7.25 34 26.5 36.975 ;
        RECT 7.2 34 26.5 36.925 ;
        RECT 7.15 34 26.5 36.875 ;
        RECT 7.1 34 26.5 36.825 ;
        RECT 7.05 34 26.5 36.775 ;
        RECT 7 34 26.5 36.725 ;
        RECT 6.95 34 26.5 36.675 ;
        RECT 6.9 34 26.5 36.625 ;
        RECT 6.85 34 26.5 36.575 ;
        RECT 6.8 34 26.5 36.525 ;
        RECT 6.75 34 26.5 36.475 ;
        RECT 6.7 34 26.5 36.425 ;
        RECT 6.65 34 26.5 36.375 ;
        RECT 6.6 34 26.5 36.325 ;
        RECT 6.55 34 26.5 36.275 ;
        RECT 6.5 34 26.5 36.225 ;
        RECT 6.45 34 26.5 36.175 ;
        RECT 6.4 34 26.5 36.125 ;
        RECT 6.35 34 26.5 36.075 ;
        RECT 6.3 34 26.5 36.025 ;
        RECT 6.25 34 26.5 35.975 ;
        RECT 6.2 34 26.5 35.925 ;
        RECT 6.15 34 26.5 35.875 ;
        RECT 6.1 34 26.5 35.825 ;
        RECT 6.05 34 26.5 35.775 ;
        RECT 6 34 26.5 35.725 ;
        RECT 5.95 34 26.5 35.675 ;
        RECT 5.9 34 26.5 35.625 ;
        RECT 5.85 34 26.5 35.575 ;
        RECT 5.8 34 26.5 35.525 ;
        RECT 5.75 34 26.5 35.475 ;
        RECT 5.7 34 26.5 35.425 ;
        RECT 5.65 34 26.5 35.375 ;
        RECT 5.6 34 26.5 35.325 ;
        RECT 5.55 34 26.5 35.275 ;
        RECT 5.5 34 26.5 35.225 ;
        RECT 1.3 0 5.5 31.025 ;
        RECT 5.45 34 26.5 35.175 ;
        RECT 5.4 34 26.5 35.125 ;
        RECT 5.35 34 26.5 35.075 ;
        RECT 5.3 34 26.5 35.025 ;
        RECT 5.25 34 26.5 34.975 ;
        RECT 5.2 34 26.5 34.925 ;
        RECT 5.15 34 26.5 34.875 ;
        RECT 5.1 34 26.5 34.825 ;
        RECT 5.05 34 26.5 34.775 ;
        RECT 5 34 26.5 34.725 ;
        RECT 4.95 34 26.5 34.675 ;
        RECT 4.9 34 26.5 34.625 ;
        RECT 4.85 34 26.5 34.575 ;
        RECT 4.8 34 26.5 34.525 ;
        RECT 4.75 34 26.5 34.475 ;
        RECT 4.7 34 26.5 34.425 ;
        RECT 4.65 34 26.5 34.375 ;
        RECT 4.6 34 26.5 34.325 ;
        RECT 4.55 34 26.5 34.275 ;
        RECT 4.5 34 26.5 34.225 ;
        RECT 4.45 34 26.5 34.175 ;
        RECT 4.4 34 26.5 34.125 ;
        RECT 4.35 34 26.5 34.075 ;
        RECT 4.25 27 12.5 33.975 ;
        RECT 4.2 27 12.5 33.925 ;
        RECT 4.15 27 12.5 33.875 ;
        RECT 4.1 27 12.5 33.825 ;
        RECT 4.05 27 12.5 33.775 ;
        RECT 4 27 12.5 33.725 ;
        RECT 3.95 27 12.5 33.675 ;
        RECT 3.9 27 12.5 33.625 ;
        RECT 3.85 27 12.5 33.575 ;
        RECT 3.8 27 12.5 33.525 ;
        RECT 3.75 27 12.5 33.475 ;
        RECT 3.7 27 12.5 33.425 ;
        RECT 3.65 27 12.5 33.375 ;
        RECT 3.6 27 12.5 33.325 ;
        RECT 3.55 27 12.5 33.275 ;
        RECT 3.5 27 12.5 33.225 ;
        RECT 3.45 27 12.5 33.175 ;
        RECT 3.4 27 12.5 33.125 ;
        RECT 3.35 27 12.5 33.075 ;
        RECT 3.3 27 12.5 33.025 ;
        RECT 3.25 27 12.5 32.975 ;
        RECT 3.2 27 12.5 32.925 ;
        RECT 3.15 27 12.5 32.875 ;
        RECT 3.1 27 12.5 32.825 ;
        RECT 3.05 27 12.5 32.775 ;
        RECT 3 27 12.5 32.725 ;
        RECT 2.95 27 12.5 32.675 ;
        RECT 2.9 27 12.5 32.625 ;
        RECT 2.85 27 12.5 32.575 ;
        RECT 2.8 27 12.5 32.525 ;
        RECT 2.75 27 12.5 32.475 ;
        RECT 2.7 27 12.5 32.425 ;
        RECT 2.65 27 12.5 32.375 ;
        RECT 2.6 27 12.5 32.325 ;
        RECT 2.55 27 12.5 32.275 ;
        RECT 2.5 27 12.5 32.225 ;
        RECT 2.45 27 12.5 32.175 ;
        RECT 2.4 27 12.5 32.125 ;
        RECT 2.35 27 12.5 32.075 ;
        RECT 2.3 27 12.5 32.025 ;
        RECT 2.25 27 12.5 31.975 ;
        RECT 2.2 27 12.5 31.925 ;
        RECT 2.15 27 12.5 31.875 ;
        RECT 2.1 27 12.5 31.825 ;
        RECT 2.05 27 12.5 31.775 ;
        RECT 2 27 12.5 31.725 ;
        RECT 1.95 27 12.5 31.675 ;
        RECT 1.9 27 12.5 31.625 ;
        RECT 1.85 27 12.5 31.575 ;
        RECT 1.8 27 12.5 31.525 ;
        RECT 1.75 27 12.5 31.475 ;
        RECT 1.7 27 12.5 31.425 ;
        RECT 1.65 27 12.5 31.375 ;
        RECT 1.6 27 12.5 31.325 ;
        RECT 1.55 27 12.5 31.275 ;
        RECT 1.5 27 12.5 31.225 ;
        RECT 1.45 27 12.5 31.175 ;
        RECT 1.4 27 12.5 31.125 ;
        RECT 1.35 27 12.5 31.075 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 29 0 48 2.5 ;
        RECT 47.5 0 48 28.5 ;
        RECT 29 0 75.5 0.5 ;
    END
  END gnd
  OBS
    LAYER M1 ;
      RECT 1.3 0 48 74.7 ;
    LAYER M2 ;
      RECT 1.3 0 48 74.7 ;
    LAYER M3 ;
      RECT 1.3 0 48 74.7 ;
    LAYER M4 ;
      RECT 1.3 0 48 74.7 ;
    LAYER M5 ;
      RECT 1.3 0 48 74.7 ;
    LAYER M6 ;
      RECT 1.3 0 48 74.7 ;
    LAYER M7 ;
      RECT 1.3 0 48 74.7 ;
    LAYER AP ;
      RECT 1.3 0 48 74.7 ;
  END
END PADSPACE_C_74x48u_CH_Rot

MACRO PADSPACE_74x6u
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN PADSPACE_74x6u 0 0 ;
  SIZE 6 BY 74 ;
  SYMMETRY X Y R90 ;
  SITE IOSite ;
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 0 1.3 1.065 26.5 ;
        RECT 5 1.3 6 26.5 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 0 29 1 74 ;
        RECT 5 29 6 74 ;
    END
  END gnd
  OBS
    LAYER M1 ;
      RECT 0 0 6 74 ;
    LAYER M2 ;
      RECT 0 0 6 74 ;
    LAYER M3 ;
      RECT 0 0 6 74 ;
    LAYER M4 ;
      RECT 0 0 6 74 ;
    LAYER M5 ;
      RECT 0 0 6 74 ;
    LAYER M6 ;
      RECT 0 0 6 74 ;
    LAYER M7 ;
      RECT 0 0 6 74 ;
    LAYER AP ;
      RECT 0 0 6 74 ;
  END
END PADSPACE_74x6u

MACRO PADSPACE_74x8u
    CLASS PAD SPACER ;
    FOREIGN PADSPACE_74x8u 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.000 BY 74.200 ;
    SYMMETRY R90 ;
    SITE IOSite ;
    PIN gnd
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M1 ;
        RECT  7.500 29.000 8.000 75.500 ;
        RECT  6.000 29.000 8.000 45.910 ;
        RECT  0.000 29.000 2.000 45.910 ;
        RECT  0.000 71.590 1.500 72.410 ;
        RECT  0.000 64.590 1.500 65.410 ;
        RECT  0.000 57.590 1.500 58.410 ;
        RECT  0.000 50.590 1.500 51.410 ;
        RECT  0.000 29.000 0.500 75.500 ;
        END
    END gnd
    PIN vdd
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M1 ;
        RECT  7.500 1.300 8.000 26.500 ;
        RECT  0.000 22.590 1.500 23.410 ;
        RECT  0.000 15.590 1.500 16.410 ;
        RECT  0.000 8.590 1.500 9.410 ;
        RECT  0.000 1.300 0.500 26.500 ;
        END
    END vdd
    OBS
        LAYER M1 ;
        RECT  2.090 1.300 5.910 7.000 ;
        RECT  2.090 11.000 5.910 14.000 ;
        RECT  2.090 18.000 5.910 21.000 ;
        RECT  3.090 1.300 5.910 27.410 ;
        RECT  2.090 25.000 5.910 27.410 ;
        RECT  3.590 1.300 4.410 75.500 ;
        RECT  2.090 47.500 5.910 49.000 ;
        RECT  2.090 53.000 5.910 56.000 ;
        RECT  2.090 60.000 5.910 63.000 ;
        RECT  2.090 67.000 5.910 70.000 ;
        RECT  3.090 47.500 5.910 75.500 ;
        RECT  2.090 74.000 5.910 75.500 ;
        LAYER M2 ;
        RECT  0.000 1.300 8.000 26.500 ;
        RECT  1.500 1.300 6.500 28.810 ;
        RECT  0.000 36.500 8.000 37.500 ;
        RECT  0.000 39.500 8.000 40.500 ;
        RECT  2.190 1.300 5.810 75.500 ;
        RECT  1.500 46.100 6.500 75.500 ;
        RECT  0.000 47.500 8.000 75.500 ;
        LAYER M3 ;
        RECT  1.500 2.800 6.500 74.000 ;
        LAYER M4 ;
        RECT  1.500 2.800 6.500 74.000 ;
        LAYER M5 ;
        RECT  1.500 2.800 6.500 74.000 ;
        LAYER M6 ;
        RECT  1.500 2.800 6.500 74.000 ;
        LAYER M7 ;
        RECT  1.500 2.800 6.500 74.000 ;
        LAYER AP ;
        RECT  1.000 2.300 7.000 74.500 ;
    END
END PADSPACE_74x8u

MACRO PADSPACE_74x4u
    CLASS PAD SPACER ;
    FOREIGN PADSPACE_74x4u 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 74.200 ;
    SYMMETRY R90 ;
    SITE IOSite ;
    PIN gnd
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M1 ;
        RECT  3.500 29.000 4.000 75.500 ;
        RECT  0.000 29.000 0.500 75.500 ;
        END
    END gnd
    PIN vdd
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M1 ;
        RECT  3.500 1.300 4.000 26.500 ;
        RECT  0.000 1.300 0.500 26.500 ;
        END
    END vdd
    OBS
        LAYER M2 ;
        RECT  0.000 1.300 4.000 26.500 ;
        RECT  0.000 36.500 4.000 37.500 ;
        RECT  0.000 39.500 4.000 40.500 ;
        RECT  1.500 1.300 2.500 75.500 ;
        RECT  0.000 47.500 4.000 75.500 ;
        LAYER M3 ;
        RECT  1.500 2.800 2.500 74.000 ;
        LAYER M4 ;
        RECT  1.500 2.800 2.500 74.000 ;
        LAYER M5 ;
        RECT  1.500 2.800 2.500 74.000 ;
        LAYER M6 ;
        RECT  1.500 2.800 2.500 74.000 ;
        LAYER M7 ;
        RECT  1.500 2.800 2.500 74.000 ;
        LAYER AP ;
        RECT  1.000 2.300 3.000 74.500 ;
    END
END PADSPACE_74x4u

MACRO PADSPACE_74x2u
    CLASS PAD SPACER ;
    FOREIGN PADSPACE_74x2u 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 74.200 ;
    SYMMETRY R90 ;
    SITE IOSite ;
    PIN gnd
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M1 ;
        RECT  0.000 29.000 2.000 75.500 ;
        END
    END gnd
    PIN vdd
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.300 2.000 26.500 ;
        END
    END vdd
    OBS
        LAYER M2 ;
        RECT  0.000 47.500 2.000 75.500 ;
        RECT  0.000 39.500 2.000 40.500 ;
        RECT  0.000 36.500 2.000 37.500 ;
        RECT  0.000 1.300 2.000 26.500 ;
    END
END PADSPACE_74x2u

MACRO PADSPACE_74x1u
    CLASS PAD SPACER ;
    FOREIGN PADSPACE_74x1u 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.000 BY 74.200 ;
    SYMMETRY R90 ;
    SITE IOSite ;
    PIN gnd
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M1 ;
        RECT  0.000 29.000 1.000 75.500 ;
        END
    END gnd
    PIN vdd
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M1 ;
        RECT  0.000 1.300 1.000 26.500 ;
        END
    END vdd
    OBS
        LAYER M2 ;
        RECT  0.000 47.500 1.000 75.500 ;
        RECT  0.000 39.500 1.000 40.500 ;
        RECT  0.000 36.500 1.000 37.500 ;
        RECT  0.000 1.300 1.000 26.500 ;
    END
END PADSPACE_74x1u

MACRO PADSPACE_74x16u
    CLASS PAD SPACER ;
    FOREIGN PADSPACE_74x16u 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.000 BY 74.200 ;
    SYMMETRY R90 ;
    SITE IOSite ;
    PIN gnd
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M1 ;
        RECT  15.500 29.000 16.000 75.500 ;
        RECT  14.500 71.590 16.000 72.410 ;
        RECT  14.500 64.590 16.000 65.410 ;
        RECT  14.500 57.590 16.000 58.410 ;
        RECT  14.500 50.590 16.000 51.410 ;
        RECT  14.000 29.000 16.000 45.910 ;
        RECT  0.000 29.000 0.500 75.500 ;
        END
    END gnd
    PIN vdd
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M1 ;
        RECT  15.500 1.300 16.000 26.500 ;
        RECT  14.500 22.590 16.000 23.410 ;
        RECT  14.500 15.590 16.000 16.410 ;
        RECT  14.500 8.590 16.000 9.410 ;
        RECT  0.000 1.300 0.500 26.500 ;
        END
    END vdd
    OBS
        LAYER M1 ;
        RECT  2.090 1.300 13.910 7.000 ;
        RECT  2.090 11.000 13.910 14.000 ;
        RECT  2.090 18.000 13.910 21.000 ;
        RECT  2.090 1.300 12.910 27.410 ;
        RECT  2.090 25.000 13.910 27.410 ;
        RECT  2.090 1.300 12.410 75.500 ;
        RECT  2.090 47.500 13.910 49.000 ;
        RECT  2.090 53.000 13.910 56.000 ;
        RECT  2.090 60.000 13.910 63.000 ;
        RECT  2.090 67.000 13.910 70.000 ;
        RECT  2.090 47.500 12.910 75.500 ;
        RECT  2.090 74.000 13.910 75.500 ;
        LAYER M2 ;
        RECT  0.000 1.300 16.000 26.500 ;
        RECT  1.500 1.300 14.500 28.810 ;
        RECT  0.000 36.500 16.000 37.500 ;
        RECT  0.000 39.500 16.000 40.500 ;
        RECT  1.500 1.300 13.810 75.500 ;
        RECT  1.500 46.100 14.500 75.500 ;
        RECT  0.000 47.500 16.000 75.500 ;
        LAYER M3 ;
        RECT  1.500 2.800 14.500 74.000 ;
        LAYER M4 ;
        RECT  1.500 2.800 14.500 74.000 ;
        LAYER M5 ;
        RECT  1.500 2.800 14.500 74.000 ;
        LAYER M6 ;
        RECT  1.500 2.800 14.500 74.000 ;
        LAYER M7 ;
        RECT  1.500 2.800 14.500 74.000 ;
        LAYER AP ;
        RECT  1.000 2.300 15.000 74.500 ;
    END
END PADSPACE_74x16u

MACRO PADGND_74x50uNOTRIG
    CLASS PAD ;
    FOREIGN PADGND_74x50uNOTRIG 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 60.000 BY 75.500 ;
    SYMMETRY R90 ;
    SITE IOSite ;
    PIN gnd
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M1 ;
        RECT  59.495 29.000 60.000 75.500 ;
        RECT  0.000 29.000 0.500 75.500 ;
        END
    END gnd
    PIN GNDC
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
            CLASS CORE ;
        LAYER AP ;
        RECT  32.445 71.000 55.000 74.000 ;
        RECT  5.000 71.000 27.475 74.000 ;
        END
        PORT
            CLASS CORE ;
        LAYER M7 ;
        RECT  31.000 69.665 53.000 72.000 ;
        RECT  7.000 69.665 29.000 72.000 ;
        END
    END GNDC
    PIN vdd
        DIRECTION INOUT ;
        USE POWER ;
        PORT
            CLASS CORE ;
        LAYER M1 ;
        RECT  59.500 1.300 60.000 26.500 ;
        RECT  0.000 1.300 0.500 26.500 ;
        END
    END vdd
    OBS
        LAYER M1 ;
        RECT  2.090 1.300 57.910 27.410 ;
        RECT  2.090 1.300 57.905 75.500 ;
        LAYER M2 ;
        RECT  0.000 1.300 60.000 26.500 ;
        RECT  0.000 36.500 60.000 37.500 ;
        RECT  0.000 39.500 60.000 40.500 ;
        RECT  1.500 1.300 58.500 75.500 ;
        RECT  0.000 47.500 60.000 75.500 ;
        LAYER M3 ;
        RECT  1.500 1.500 58.500 74.000 ;
        LAYER M4 ;
        RECT  1.500 1.500 58.500 74.000 ;
        LAYER M5 ;
        RECT  1.500 1.500 58.500 74.000 ;
        RECT  2.000 1.500 58.000 75.500 ;
        LAYER M6 ;
        RECT  1.500 1.500 58.500 74.000 ;
        RECT  2.000 1.500 58.000 75.500 ;
        LAYER M7 ;
        RECT  5.500 1.300 47.500 65.965 ;
        RECT  1.500 1.500 58.500 65.965 ;
        RECT  1.500 1.500 3.300 74.000 ;
        RECT  56.700 1.500 58.500 74.000 ;
        LAYER AP ;
        RECT  1.000 1.000 59.000 65.465 ;
        RECT  1.000 1.000 2.800 66.800 ;
        RECT  5.000 0.000 55.000 66.800 ;
        RECT  57.200 1.000 59.000 66.800 ;
    END
END PADGND_74x50uNOTRIG

MACRO CPAD_S_74x50u_GND
    CLASS PAD ;
    FOREIGN CPAD_S_74x50u_VDD 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 50.000 BY 75.500 ;
    SYMMETRY R90 ;
    SITE IOSite ;
    PIN gnd
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M1 ;
        RECT  49.500 29.000 50.000 75.500 ;
        RECT  48.000 71.590 50.000 72.410 ;
        RECT  48.000 64.590 50.000 65.410 ;
        RECT  48.000 57.590 50.000 58.410 ;
        RECT  48.000 50.590 50.000 51.410 ;
        RECT  0.000 71.590 2.000 72.410 ;
        RECT  0.000 64.590 2.000 65.410 ;
        RECT  0.000 57.590 2.000 58.410 ;
        RECT  0.000 50.590 2.000 51.410 ;
        RECT  0.000 29.000 2.000 45.910 ;
        RECT  0.000 29.000 0.500 75.500 ;
        END
    END gnd
    PIN vdd
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M1 ;
        RECT  49.500 1.300 50.000 26.500 ;
        RECT  48.000 22.590 50.000 23.410 ;
        RECT  48.000 15.590 50.000 16.410 ;
        RECT  48.000 8.590 50.000 9.410 ;
        RECT  0.000 22.590 2.000 23.410 ;
        RECT  0.000 15.590 2.000 16.410 ;
        RECT  0.000 8.590 2.000 9.410 ;
        RECT  0.000 1.300 0.500 26.500 ;
        END
    END vdd
    PIN GNDC
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
            CLASS CORE ;
        LAYER AP ;
        RECT  27.480 71.000 50.000 74.000 ;
        RECT  0.000 71.000 22.510 74.000 ;
        END
        PORT
            CLASS CORE ;
        LAYER M7 ;
        RECT  26.000 69.665 48.000 72.000 ;
        RECT  2.000 69.665 24.000 72.000 ;
        END
    END GNDC
    OBS
        LAYER M1 ;
        RECT  2.090 1.300 47.910 7.000 ;
        RECT  2.090 11.000 47.910 14.000 ;
        RECT  2.090 18.000 47.910 21.000 ;
        RECT  2.090 25.000 47.910 27.410 ;
        RECT  3.590 25.000 47.910 49.000 ;
        RECT  2.090 47.500 47.910 49.000 ;
        RECT  2.090 53.000 47.910 56.000 ;
        RECT  2.090 60.000 47.910 63.000 ;
        RECT  2.090 67.000 47.910 70.000 ;
        RECT  3.590 1.300 46.410 75.500 ;
        RECT  2.090 74.000 47.910 75.500 ;
        LAYER M2 ;
        RECT  0.000 1.300 50.000 26.500 ;
        RECT  1.500 1.300 48.500 28.810 ;
        RECT  0.000 36.500 50.000 37.500 ;
        RECT  0.000 39.500 50.000 40.500 ;
        RECT  2.190 1.300 48.500 75.500 ;
        RECT  1.500 46.100 48.500 75.500 ;
        RECT  0.000 47.500 50.000 75.500 ;
        LAYER M3 ;
        RECT  1.500 1.500 48.500 74.000 ;
        LAYER M4 ;
        RECT  1.500 1.500 48.500 74.000 ;
        LAYER M5 ;
        RECT  1.500 1.500 48.500 74.000 ;
        LAYER M6 ;
        RECT  1.500 1.500 48.500 74.000 ;
        LAYER M7 ;
        RECT  3.000 1.300 42.500 65.965 ;
        RECT  1.500 1.500 48.500 65.965 ;
        RECT  0.500 5.500 49.500 65.965 ;
        LAYER AP ;
        RECT  0.000 0.000 50.000 66.800 ;
    END
END CPAD_S_74x50u_GND

MACRO CPAD_S_74x50u_VDD
    CLASS PAD ;
    FOREIGN CPAD_S_74x50u_VDD 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 50.000 BY 75.500 ;
    SYMMETRY R90 ;
    SITE IOSite ;
    PIN gnd
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M1 ;
        RECT  49.500 29.000 50.000 75.500 ;
        RECT  48.000 71.590 50.000 72.410 ;
        RECT  48.000 64.590 50.000 65.410 ;
        RECT  48.000 57.590 50.000 58.410 ;
        RECT  48.000 50.590 50.000 51.410 ;
        RECT  0.000 71.590 2.000 72.410 ;
        RECT  0.000 64.590 2.000 65.410 ;
        RECT  0.000 57.590 2.000 58.410 ;
        RECT  0.000 50.590 2.000 51.410 ;
        RECT  0.000 29.000 2.000 45.910 ;
        RECT  0.000 29.000 0.500 75.500 ;
        END
    END gnd
    PIN vdd
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M1 ;
        RECT  49.500 1.300 50.000 26.500 ;
        RECT  48.000 22.590 50.000 23.410 ;
        RECT  48.000 15.590 50.000 16.410 ;
        RECT  48.000 8.590 50.000 9.410 ;
        RECT  0.000 22.590 2.000 23.410 ;
        RECT  0.000 15.590 2.000 16.410 ;
        RECT  0.000 8.590 2.000 9.410 ;
        RECT  0.000 1.300 0.500 26.500 ;
        END
    END vdd
    PIN VDDC
        DIRECTION INOUT ;
        USE POWER ;
        PORT
            CLASS CORE ;
        LAYER AP ;
        RECT  27.480 71.000 50.000 74.000 ;
        RECT  0.000 71.000 22.510 74.000 ;
        END
        PORT
            CLASS CORE ;
        LAYER M7 ;
        RECT  26.000 69.665 48.000 72.000 ;
        RECT  2.000 69.665 24.000 72.000 ;
        END
    END VDDC
    OBS
        LAYER M1 ;
        RECT  2.090 1.300 47.910 7.000 ;
        RECT  2.090 11.000 47.910 14.000 ;
        RECT  2.090 18.000 47.910 21.000 ;
        RECT  2.090 25.000 47.910 27.410 ;
        RECT  3.590 25.000 47.910 49.000 ;
        RECT  2.090 47.500 47.910 49.000 ;
        RECT  2.090 53.000 47.910 56.000 ;
        RECT  2.090 60.000 47.910 63.000 ;
        RECT  2.090 67.000 47.910 70.000 ;
        RECT  3.590 1.300 46.410 75.500 ;
        RECT  2.090 74.000 47.910 75.500 ;
        LAYER M2 ;
        RECT  0.000 1.300 50.000 26.500 ;
        RECT  1.500 1.300 48.500 28.810 ;
        RECT  0.000 36.500 50.000 37.500 ;
        RECT  0.000 39.500 50.000 40.500 ;
        RECT  2.190 1.300 48.500 75.500 ;
        RECT  1.500 46.100 48.500 75.500 ;
        RECT  0.000 47.500 50.000 75.500 ;
        LAYER M3 ;
        RECT  1.500 1.500 48.500 74.000 ;
        LAYER M4 ;
        RECT  1.500 1.500 48.500 74.000 ;
        LAYER M5 ;
        RECT  1.500 1.500 48.500 74.000 ;
        LAYER M6 ;
        RECT  1.500 1.500 48.500 74.000 ;
        LAYER M7 ;
        RECT  3.000 1.300 42.500 65.965 ;
        RECT  1.500 1.500 48.500 65.965 ;
        RECT  0.500 5.500 49.500 65.965 ;
        LAYER AP ;
        RECT  0.000 0.000 50.000 66.800 ;
    END
END CPAD_S_74x50u_VDD

MACRO CPAD_S_74x50u_OUT
    CLASS PAD ;
    FOREIGN CPAD_S_74x50u_OUT 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 50.000 BY 75.500 ;
    SYMMETRY R90 ;
    SITE IOSite ;
    PIN COREIO
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  23.090 67.675 27.090 72.000 ;
        END
    END COREIO
    PIN PADIO
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  45.795 3.300 46.500 4.045 ;
        END
    END PADIO
    PIN gnd
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M1 ;
        RECT  49.500 29.000 50.000 75.500 ;
        RECT  48.000 71.590 50.000 72.410 ;
        RECT  48.000 64.590 50.000 65.410 ;
        RECT  48.000 57.590 50.000 58.410 ;
        RECT  48.000 50.590 50.000 51.410 ;
        RECT  0.000 71.590 2.000 72.410 ;
        RECT  0.000 64.590 2.000 65.410 ;
        RECT  0.000 57.590 2.000 58.410 ;
        RECT  0.000 50.590 2.000 51.410 ;
        RECT  0.000 29.000 2.000 45.910 ;
        RECT  0.000 29.000 0.500 75.500 ;
        END
    END gnd
    PIN vdd
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M1 ;
        RECT  49.500 1.300 50.000 26.500 ;
        RECT  48.000 22.590 50.000 23.410 ;
        RECT  48.000 15.590 50.000 16.410 ;
        RECT  48.000 8.590 50.000 9.410 ;
        RECT  0.000 22.590 2.000 23.410 ;
        RECT  0.000 15.590 2.000 16.410 ;
        RECT  0.000 8.590 2.000 9.410 ;
        RECT  0.000 1.300 0.500 26.500 ;
        END
    END vdd
    OBS
        LAYER M1 ;
        RECT  2.090 1.300 47.910 7.000 ;
        RECT  2.090 11.000 47.910 14.000 ;
        RECT  2.090 18.000 47.910 21.000 ;
        RECT  2.090 25.000 47.910 27.410 ;
        RECT  3.590 25.000 47.910 49.000 ;
        RECT  2.090 47.500 47.910 49.000 ;
        RECT  2.090 53.000 47.910 56.000 ;
        RECT  2.090 60.000 47.910 63.000 ;
        RECT  2.090 67.000 47.910 70.000 ;
        RECT  3.590 1.300 46.410 75.500 ;
        RECT  2.090 74.000 47.910 75.500 ;
        LAYER M2 ;
        RECT  0.000 1.300 50.000 26.500 ;
        RECT  1.500 1.300 48.500 28.810 ;
        RECT  0.000 36.500 50.000 37.500 ;
        RECT  0.000 39.500 50.000 40.500 ;
        RECT  2.190 1.300 48.500 75.500 ;
        RECT  1.500 46.100 48.500 75.500 ;
        RECT  0.000 47.500 50.000 75.500 ;
        LAYER M3 ;
        RECT  1.500 1.500 48.500 74.000 ;
        LAYER M4 ;
        RECT  1.500 1.500 48.500 74.000 ;
        LAYER M5 ;
        RECT  1.500 1.500 48.500 74.000 ;
        LAYER M6 ;
        RECT  1.500 1.500 48.500 74.000 ;
        LAYER M7 ;
        RECT  3.000 1.300 42.095 63.975 ;
        RECT  0.500 5.500 19.390 68.500 ;
        RECT  30.790 7.745 49.500 68.500 ;
        RECT  1.500 1.500 19.390 74.000 ;
        RECT  30.790 7.745 48.500 74.000 ;
        LAYER AP ;
        RECT  0.000 0.000 50.000 74.000 ;
        RECT  1.000 0.000 18.890 74.500 ;
        RECT  31.290 0.000 49.000 74.500 ;
    END
END CPAD_S_74x50u_OUT

MACRO CPAD_S_74x50u_IN
    CLASS PAD ;
    FOREIGN CPAD_S_74x50u_IN 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 50.000 BY 75.500 ;
    SYMMETRY R90 ;
    SITE IOSite ;
    PIN COREIO
        DIRECTION OUTPUT ;
        PORT
        LAYER M7 ;
        RECT  23.075 67.540 27.075 72.000 ;
        END
    END COREIO
    PIN PADIO
        DIRECTION INPUT ;
        PORT
        LAYER M7 ;
        RECT  45.770 3.300 46.500 3.910 ;
        END
    END PADIO
    PIN gnd
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER M1 ;
        RECT  49.500 29.000 50.000 75.500 ;
        RECT  48.000 71.590 50.000 72.410 ;
        RECT  48.000 64.590 50.000 65.410 ;
        RECT  48.000 57.590 50.000 58.410 ;
        RECT  48.000 50.590 50.000 51.410 ;
        RECT  0.000 71.590 2.000 72.410 ;
        RECT  0.000 64.590 2.000 65.410 ;
        RECT  0.000 57.590 2.000 58.410 ;
        RECT  0.000 50.590 2.000 51.410 ;
        RECT  0.000 29.000 2.000 45.910 ;
        RECT  0.000 29.000 0.500 75.500 ;
        END
    END gnd
    PIN vdd
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER M1 ;
        RECT  49.500 1.300 50.000 26.500 ;
        RECT  48.000 22.590 50.000 23.410 ;
        RECT  48.000 15.590 50.000 16.410 ;
        RECT  48.000 8.590 50.000 9.410 ;
        RECT  0.000 22.590 2.000 23.410 ;
        RECT  0.000 15.590 2.000 16.410 ;
        RECT  0.000 8.590 2.000 9.410 ;
        RECT  0.000 1.300 0.500 26.500 ;
        END
    END vdd
    OBS
        LAYER M1 ;
        RECT  2.090 1.300 47.910 7.000 ;
        RECT  2.090 11.000 47.910 14.000 ;
        RECT  2.090 18.000 47.910 21.000 ;
        RECT  2.090 25.000 47.910 27.410 ;
        RECT  3.590 25.000 47.910 49.000 ;
        RECT  2.090 47.500 47.910 49.000 ;
        RECT  2.090 53.000 47.910 56.000 ;
        RECT  2.090 60.000 47.910 63.000 ;
        RECT  2.090 67.000 47.910 70.000 ;
        RECT  3.590 1.300 46.410 75.500 ;
        RECT  2.090 74.000 47.910 75.500 ;
        LAYER M2 ;
        RECT  0.000 1.300 50.000 26.500 ;
        RECT  1.500 1.300 48.500 28.810 ;
        RECT  0.000 36.500 50.000 37.500 ;
        RECT  0.000 39.500 50.000 40.500 ;
        RECT  2.190 1.300 48.500 75.500 ;
        RECT  1.500 46.100 48.500 75.500 ;
        RECT  0.000 47.500 50.000 75.500 ;
        LAYER M3 ;
        RECT  1.500 1.500 48.500 74.000 ;
        LAYER M4 ;
        RECT  1.500 1.500 48.500 74.000 ;
        LAYER M5 ;
        RECT  1.500 1.500 48.500 74.000 ;
        LAYER M6 ;
        RECT  1.500 1.500 48.500 74.000 ;
        LAYER M7 ;
        RECT  3.000 1.300 42.070 63.840 ;
        RECT  0.500 5.500 19.375 68.500 ;
        RECT  30.775 7.610 49.500 68.500 ;
        RECT  1.500 1.500 19.375 74.000 ;
        RECT  30.775 7.610 48.500 74.000 ;
        LAYER AP ;
        RECT  0.000 0.000 50.000 74.000 ;
        RECT  1.000 0.000 18.875 74.500 ;
        RECT  31.275 0.000 49.000 74.500 ;
    END
END CPAD_S_74x50u_IN

END LIBRARY
